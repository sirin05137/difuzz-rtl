module RocketTile(
  input         clock,
  input         reset,
  input         auto_intsink_in_sync_0,
  input         auto_int_in_xing_in_2_sync_0,
  input         auto_int_in_xing_in_1_sync_0,
  input         auto_int_in_xing_in_0_sync_0,
  input         auto_int_in_xing_in_0_sync_1,
  input         auto_tl_master_xing_out_a_ready,
  output        auto_tl_master_xing_out_a_valid,
  output [2:0]  auto_tl_master_xing_out_a_bits_opcode,
  output [2:0]  auto_tl_master_xing_out_a_bits_param,
  output [3:0]  auto_tl_master_xing_out_a_bits_size,
  output [1:0]  auto_tl_master_xing_out_a_bits_source,
  output [31:0] auto_tl_master_xing_out_a_bits_address,
  output [7:0]  auto_tl_master_xing_out_a_bits_mask,
  output [63:0] auto_tl_master_xing_out_a_bits_data,
  output        auto_tl_master_xing_out_a_bits_corrupt,
  output        auto_tl_master_xing_out_b_ready,
  input         auto_tl_master_xing_out_b_valid,
  input  [2:0]  auto_tl_master_xing_out_b_bits_opcode,
  input  [1:0]  auto_tl_master_xing_out_b_bits_param,
  input  [3:0]  auto_tl_master_xing_out_b_bits_size,
  input  [1:0]  auto_tl_master_xing_out_b_bits_source,
  input  [31:0] auto_tl_master_xing_out_b_bits_address,
  input  [7:0]  auto_tl_master_xing_out_b_bits_mask,
  input  [63:0] auto_tl_master_xing_out_b_bits_data,
  input         auto_tl_master_xing_out_b_bits_corrupt,
  input         auto_tl_master_xing_out_c_ready,
  output        auto_tl_master_xing_out_c_valid,
  output [2:0]  auto_tl_master_xing_out_c_bits_opcode,
  output [2:0]  auto_tl_master_xing_out_c_bits_param,
  output [3:0]  auto_tl_master_xing_out_c_bits_size,
  output [1:0]  auto_tl_master_xing_out_c_bits_source,
  output [31:0] auto_tl_master_xing_out_c_bits_address,
  output [63:0] auto_tl_master_xing_out_c_bits_data,
  output        auto_tl_master_xing_out_c_bits_corrupt,
  output        auto_tl_master_xing_out_d_ready,
  input         auto_tl_master_xing_out_d_valid,
  input  [2:0]  auto_tl_master_xing_out_d_bits_opcode,
  input  [1:0]  auto_tl_master_xing_out_d_bits_param,
  input  [3:0]  auto_tl_master_xing_out_d_bits_size,
  input  [1:0]  auto_tl_master_xing_out_d_bits_source,
  input  [1:0]  auto_tl_master_xing_out_d_bits_sink,
  input         auto_tl_master_xing_out_d_bits_denied,
  input  [63:0] auto_tl_master_xing_out_d_bits_data,
  input         auto_tl_master_xing_out_d_bits_corrupt,
  input         auto_tl_master_xing_out_e_ready,
  output        auto_tl_master_xing_out_e_valid,
  output [1:0]  auto_tl_master_xing_out_e_bits_sink,
  input  [1:0]  constants_hartid,
  input  [31:0] constants_reset_vector,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         intsink_1_halt,
  input         intsink_halt,
  input         dcache_halt,
  input         dcacheArb_halt,
  input         intsink_2_halt,
  input         frontend_halt,
  input         buffer_halt,
  input         core_halt,
  input         intsink_3_halt,
  input         ptw_halt,
  input         tlMasterXbar_halt,
  input         fpuOpt_halt,
  input         intXbar_halt
);
  wire  tlMasterXbar_clock; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_reset; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_in_1_a_ready; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_in_1_a_valid; // @[BaseTile.scala 142:42]
  wire [31:0] tlMasterXbar_auto_in_1_a_bits_address; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_in_1_d_valid; // @[BaseTile.scala 142:42]
  wire [2:0] tlMasterXbar_auto_in_1_d_bits_opcode; // @[BaseTile.scala 142:42]
  wire [3:0] tlMasterXbar_auto_in_1_d_bits_size; // @[BaseTile.scala 142:42]
  wire [63:0] tlMasterXbar_auto_in_1_d_bits_data; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_in_1_d_bits_corrupt; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_in_0_a_ready; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_in_0_a_valid; // @[BaseTile.scala 142:42]
  wire [2:0] tlMasterXbar_auto_in_0_a_bits_opcode; // @[BaseTile.scala 142:42]
  wire [2:0] tlMasterXbar_auto_in_0_a_bits_param; // @[BaseTile.scala 142:42]
  wire [3:0] tlMasterXbar_auto_in_0_a_bits_size; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_in_0_a_bits_source; // @[BaseTile.scala 142:42]
  wire [31:0] tlMasterXbar_auto_in_0_a_bits_address; // @[BaseTile.scala 142:42]
  wire [7:0] tlMasterXbar_auto_in_0_a_bits_mask; // @[BaseTile.scala 142:42]
  wire [63:0] tlMasterXbar_auto_in_0_a_bits_data; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_in_0_b_ready; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_in_0_b_valid; // @[BaseTile.scala 142:42]
  wire [1:0] tlMasterXbar_auto_in_0_b_bits_param; // @[BaseTile.scala 142:42]
  wire [3:0] tlMasterXbar_auto_in_0_b_bits_size; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_in_0_b_bits_source; // @[BaseTile.scala 142:42]
  wire [31:0] tlMasterXbar_auto_in_0_b_bits_address; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_in_0_c_ready; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_in_0_c_valid; // @[BaseTile.scala 142:42]
  wire [2:0] tlMasterXbar_auto_in_0_c_bits_opcode; // @[BaseTile.scala 142:42]
  wire [2:0] tlMasterXbar_auto_in_0_c_bits_param; // @[BaseTile.scala 142:42]
  wire [3:0] tlMasterXbar_auto_in_0_c_bits_size; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_in_0_c_bits_source; // @[BaseTile.scala 142:42]
  wire [31:0] tlMasterXbar_auto_in_0_c_bits_address; // @[BaseTile.scala 142:42]
  wire [63:0] tlMasterXbar_auto_in_0_c_bits_data; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_in_0_d_ready; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_in_0_d_valid; // @[BaseTile.scala 142:42]
  wire [2:0] tlMasterXbar_auto_in_0_d_bits_opcode; // @[BaseTile.scala 142:42]
  wire [1:0] tlMasterXbar_auto_in_0_d_bits_param; // @[BaseTile.scala 142:42]
  wire [3:0] tlMasterXbar_auto_in_0_d_bits_size; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_in_0_d_bits_source; // @[BaseTile.scala 142:42]
  wire [1:0] tlMasterXbar_auto_in_0_d_bits_sink; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_in_0_d_bits_denied; // @[BaseTile.scala 142:42]
  wire [63:0] tlMasterXbar_auto_in_0_d_bits_data; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_in_0_e_ready; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_in_0_e_valid; // @[BaseTile.scala 142:42]
  wire [1:0] tlMasterXbar_auto_in_0_e_bits_sink; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_out_a_ready; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_out_a_valid; // @[BaseTile.scala 142:42]
  wire [2:0] tlMasterXbar_auto_out_a_bits_opcode; // @[BaseTile.scala 142:42]
  wire [2:0] tlMasterXbar_auto_out_a_bits_param; // @[BaseTile.scala 142:42]
  wire [3:0] tlMasterXbar_auto_out_a_bits_size; // @[BaseTile.scala 142:42]
  wire [1:0] tlMasterXbar_auto_out_a_bits_source; // @[BaseTile.scala 142:42]
  wire [31:0] tlMasterXbar_auto_out_a_bits_address; // @[BaseTile.scala 142:42]
  wire [7:0] tlMasterXbar_auto_out_a_bits_mask; // @[BaseTile.scala 142:42]
  wire [63:0] tlMasterXbar_auto_out_a_bits_data; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_out_a_bits_corrupt; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_out_b_ready; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_out_b_valid; // @[BaseTile.scala 142:42]
  wire [2:0] tlMasterXbar_auto_out_b_bits_opcode; // @[BaseTile.scala 142:42]
  wire [1:0] tlMasterXbar_auto_out_b_bits_param; // @[BaseTile.scala 142:42]
  wire [3:0] tlMasterXbar_auto_out_b_bits_size; // @[BaseTile.scala 142:42]
  wire [1:0] tlMasterXbar_auto_out_b_bits_source; // @[BaseTile.scala 142:42]
  wire [31:0] tlMasterXbar_auto_out_b_bits_address; // @[BaseTile.scala 142:42]
  wire [7:0] tlMasterXbar_auto_out_b_bits_mask; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_out_b_bits_corrupt; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_out_c_ready; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_out_c_valid; // @[BaseTile.scala 142:42]
  wire [2:0] tlMasterXbar_auto_out_c_bits_opcode; // @[BaseTile.scala 142:42]
  wire [2:0] tlMasterXbar_auto_out_c_bits_param; // @[BaseTile.scala 142:42]
  wire [3:0] tlMasterXbar_auto_out_c_bits_size; // @[BaseTile.scala 142:42]
  wire [1:0] tlMasterXbar_auto_out_c_bits_source; // @[BaseTile.scala 142:42]
  wire [31:0] tlMasterXbar_auto_out_c_bits_address; // @[BaseTile.scala 142:42]
  wire [63:0] tlMasterXbar_auto_out_c_bits_data; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_out_d_ready; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_out_d_valid; // @[BaseTile.scala 142:42]
  wire [2:0] tlMasterXbar_auto_out_d_bits_opcode; // @[BaseTile.scala 142:42]
  wire [1:0] tlMasterXbar_auto_out_d_bits_param; // @[BaseTile.scala 142:42]
  wire [3:0] tlMasterXbar_auto_out_d_bits_size; // @[BaseTile.scala 142:42]
  wire [1:0] tlMasterXbar_auto_out_d_bits_source; // @[BaseTile.scala 142:42]
  wire [1:0] tlMasterXbar_auto_out_d_bits_sink; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_out_d_bits_denied; // @[BaseTile.scala 142:42]
  wire [63:0] tlMasterXbar_auto_out_d_bits_data; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_out_d_bits_corrupt; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_out_e_ready; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_auto_out_e_valid; // @[BaseTile.scala 142:42]
  wire [1:0] tlMasterXbar_auto_out_e_bits_sink; // @[BaseTile.scala 142:42]
  wire [29:0] tlMasterXbar_io_covSum; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_metaAssert; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_metaReset; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_TLMonitor_halt; // @[BaseTile.scala 142:42]
  wire  tlMasterXbar_TLMonitor_1_halt; // @[BaseTile.scala 142:42]
  wire  intXbar_auto_int_in_3_0; // @[BaseTile.scala 144:37]
  wire  intXbar_auto_int_in_2_0; // @[BaseTile.scala 144:37]
  wire  intXbar_auto_int_in_1_0; // @[BaseTile.scala 144:37]
  wire  intXbar_auto_int_in_1_1; // @[BaseTile.scala 144:37]
  wire  intXbar_auto_int_in_0_0; // @[BaseTile.scala 144:37]
  wire  intXbar_auto_int_out_0; // @[BaseTile.scala 144:37]
  wire  intXbar_auto_int_out_1; // @[BaseTile.scala 144:37]
  wire  intXbar_auto_int_out_2; // @[BaseTile.scala 144:37]
  wire  intXbar_auto_int_out_3; // @[BaseTile.scala 144:37]
  wire  intXbar_auto_int_out_4; // @[BaseTile.scala 144:37]
  wire [29:0] intXbar_io_covSum; // @[BaseTile.scala 144:37]
  wire  intXbar_metaAssert; // @[BaseTile.scala 144:37]
  wire  dcache_gated_clock; // @[HellaCache.scala 215:43]
  wire  dcache_reset; // @[HellaCache.scala 215:43]
  wire  dcache_auto_out_a_ready; // @[HellaCache.scala 215:43]
  wire  dcache_auto_out_a_valid; // @[HellaCache.scala 215:43]
  wire [2:0] dcache_auto_out_a_bits_opcode; // @[HellaCache.scala 215:43]
  wire [2:0] dcache_auto_out_a_bits_param; // @[HellaCache.scala 215:43]
  wire [3:0] dcache_auto_out_a_bits_size; // @[HellaCache.scala 215:43]
  wire  dcache_auto_out_a_bits_source; // @[HellaCache.scala 215:43]
  wire [31:0] dcache_auto_out_a_bits_address; // @[HellaCache.scala 215:43]
  wire [7:0] dcache_auto_out_a_bits_mask; // @[HellaCache.scala 215:43]
  wire [63:0] dcache_auto_out_a_bits_data; // @[HellaCache.scala 215:43]
  wire  dcache_auto_out_b_ready; // @[HellaCache.scala 215:43]
  wire  dcache_auto_out_b_valid; // @[HellaCache.scala 215:43]
  wire [1:0] dcache_auto_out_b_bits_param; // @[HellaCache.scala 215:43]
  wire [3:0] dcache_auto_out_b_bits_size; // @[HellaCache.scala 215:43]
  wire  dcache_auto_out_b_bits_source; // @[HellaCache.scala 215:43]
  wire [31:0] dcache_auto_out_b_bits_address; // @[HellaCache.scala 215:43]
  wire  dcache_auto_out_c_ready; // @[HellaCache.scala 215:43]
  wire  dcache_auto_out_c_valid; // @[HellaCache.scala 215:43]
  wire [2:0] dcache_auto_out_c_bits_opcode; // @[HellaCache.scala 215:43]
  wire [2:0] dcache_auto_out_c_bits_param; // @[HellaCache.scala 215:43]
  wire [3:0] dcache_auto_out_c_bits_size; // @[HellaCache.scala 215:43]
  wire  dcache_auto_out_c_bits_source; // @[HellaCache.scala 215:43]
  wire [31:0] dcache_auto_out_c_bits_address; // @[HellaCache.scala 215:43]
  wire [63:0] dcache_auto_out_c_bits_data; // @[HellaCache.scala 215:43]
  wire  dcache_auto_out_d_ready; // @[HellaCache.scala 215:43]
  wire  dcache_auto_out_d_valid; // @[HellaCache.scala 215:43]
  wire [2:0] dcache_auto_out_d_bits_opcode; // @[HellaCache.scala 215:43]
  wire [1:0] dcache_auto_out_d_bits_param; // @[HellaCache.scala 215:43]
  wire [3:0] dcache_auto_out_d_bits_size; // @[HellaCache.scala 215:43]
  wire  dcache_auto_out_d_bits_source; // @[HellaCache.scala 215:43]
  wire [1:0] dcache_auto_out_d_bits_sink; // @[HellaCache.scala 215:43]
  wire  dcache_auto_out_d_bits_denied; // @[HellaCache.scala 215:43]
  wire [63:0] dcache_auto_out_d_bits_data; // @[HellaCache.scala 215:43]
  wire  dcache_auto_out_e_ready; // @[HellaCache.scala 215:43]
  wire  dcache_auto_out_e_valid; // @[HellaCache.scala 215:43]
  wire [1:0] dcache_auto_out_e_bits_sink; // @[HellaCache.scala 215:43]
  wire  dcache_io_cpu_req_ready; // @[HellaCache.scala 215:43]
  wire  dcache_io_cpu_req_valid; // @[HellaCache.scala 215:43]
  wire [39:0] dcache_io_cpu_req_bits_addr; // @[HellaCache.scala 215:43]
  wire [6:0] dcache_io_cpu_req_bits_tag; // @[HellaCache.scala 215:43]
  wire [4:0] dcache_io_cpu_req_bits_cmd; // @[HellaCache.scala 215:43]
  wire [2:0] dcache_io_cpu_req_bits_typ; // @[HellaCache.scala 215:43]
  wire  dcache_io_cpu_req_bits_phys; // @[HellaCache.scala 215:43]
  wire  dcache_io_cpu_s1_kill; // @[HellaCache.scala 215:43]
  wire [63:0] dcache_io_cpu_s1_data_data; // @[HellaCache.scala 215:43]
  wire  dcache_io_cpu_s2_nack; // @[HellaCache.scala 215:43]
  wire  dcache_io_cpu_resp_valid; // @[HellaCache.scala 215:43]
  wire [6:0] dcache_io_cpu_resp_bits_tag; // @[HellaCache.scala 215:43]
  wire [2:0] dcache_io_cpu_resp_bits_typ; // @[HellaCache.scala 215:43]
  wire [63:0] dcache_io_cpu_resp_bits_data; // @[HellaCache.scala 215:43]
  wire  dcache_io_cpu_resp_bits_replay; // @[HellaCache.scala 215:43]
  wire  dcache_io_cpu_resp_bits_has_data; // @[HellaCache.scala 215:43]
  wire [63:0] dcache_io_cpu_resp_bits_data_word_bypass; // @[HellaCache.scala 215:43]
  wire  dcache_io_cpu_replay_next; // @[HellaCache.scala 215:43]
  wire  dcache_io_cpu_s2_xcpt_ma_ld; // @[HellaCache.scala 215:43]
  wire  dcache_io_cpu_s2_xcpt_ma_st; // @[HellaCache.scala 215:43]
  wire  dcache_io_cpu_s2_xcpt_pf_ld; // @[HellaCache.scala 215:43]
  wire  dcache_io_cpu_s2_xcpt_pf_st; // @[HellaCache.scala 215:43]
  wire  dcache_io_cpu_s2_xcpt_ae_ld; // @[HellaCache.scala 215:43]
  wire  dcache_io_cpu_s2_xcpt_ae_st; // @[HellaCache.scala 215:43]
  wire  dcache_io_cpu_ordered; // @[HellaCache.scala 215:43]
  wire  dcache_io_cpu_perf_grant; // @[HellaCache.scala 215:43]
  wire  dcache_io_cpu_keep_clock_enabled; // @[HellaCache.scala 215:43]
  wire  dcache_io_cpu_clock_enabled; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_req_ready; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_req_valid; // @[HellaCache.scala 215:43]
  wire [26:0] dcache_io_ptw_req_bits_bits_addr; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_resp_valid; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_resp_bits_ae; // @[HellaCache.scala 215:43]
  wire [53:0] dcache_io_ptw_resp_bits_pte_ppn; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_resp_bits_pte_d; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_resp_bits_pte_a; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_resp_bits_pte_g; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_resp_bits_pte_u; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_resp_bits_pte_x; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_resp_bits_pte_w; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_resp_bits_pte_r; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_resp_bits_pte_v; // @[HellaCache.scala 215:43]
  wire [1:0] dcache_io_ptw_resp_bits_level; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_resp_bits_homogeneous; // @[HellaCache.scala 215:43]
  wire [3:0] dcache_io_ptw_ptbr_mode; // @[HellaCache.scala 215:43]
  wire [1:0] dcache_io_ptw_status_dprv; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_status_mxr; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_status_sum; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_0_cfg_l; // @[HellaCache.scala 215:43]
  wire [1:0] dcache_io_ptw_pmp_0_cfg_a; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_0_cfg_x; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_0_cfg_w; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_0_cfg_r; // @[HellaCache.scala 215:43]
  wire [29:0] dcache_io_ptw_pmp_0_addr; // @[HellaCache.scala 215:43]
  wire [31:0] dcache_io_ptw_pmp_0_mask; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_1_cfg_l; // @[HellaCache.scala 215:43]
  wire [1:0] dcache_io_ptw_pmp_1_cfg_a; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_1_cfg_x; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_1_cfg_w; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_1_cfg_r; // @[HellaCache.scala 215:43]
  wire [29:0] dcache_io_ptw_pmp_1_addr; // @[HellaCache.scala 215:43]
  wire [31:0] dcache_io_ptw_pmp_1_mask; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_2_cfg_l; // @[HellaCache.scala 215:43]
  wire [1:0] dcache_io_ptw_pmp_2_cfg_a; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_2_cfg_x; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_2_cfg_w; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_2_cfg_r; // @[HellaCache.scala 215:43]
  wire [29:0] dcache_io_ptw_pmp_2_addr; // @[HellaCache.scala 215:43]
  wire [31:0] dcache_io_ptw_pmp_2_mask; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_3_cfg_l; // @[HellaCache.scala 215:43]
  wire [1:0] dcache_io_ptw_pmp_3_cfg_a; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_3_cfg_x; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_3_cfg_w; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_3_cfg_r; // @[HellaCache.scala 215:43]
  wire [29:0] dcache_io_ptw_pmp_3_addr; // @[HellaCache.scala 215:43]
  wire [31:0] dcache_io_ptw_pmp_3_mask; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_4_cfg_l; // @[HellaCache.scala 215:43]
  wire [1:0] dcache_io_ptw_pmp_4_cfg_a; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_4_cfg_x; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_4_cfg_w; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_4_cfg_r; // @[HellaCache.scala 215:43]
  wire [29:0] dcache_io_ptw_pmp_4_addr; // @[HellaCache.scala 215:43]
  wire [31:0] dcache_io_ptw_pmp_4_mask; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_5_cfg_l; // @[HellaCache.scala 215:43]
  wire [1:0] dcache_io_ptw_pmp_5_cfg_a; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_5_cfg_x; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_5_cfg_w; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_5_cfg_r; // @[HellaCache.scala 215:43]
  wire [29:0] dcache_io_ptw_pmp_5_addr; // @[HellaCache.scala 215:43]
  wire [31:0] dcache_io_ptw_pmp_5_mask; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_6_cfg_l; // @[HellaCache.scala 215:43]
  wire [1:0] dcache_io_ptw_pmp_6_cfg_a; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_6_cfg_x; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_6_cfg_w; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_6_cfg_r; // @[HellaCache.scala 215:43]
  wire [29:0] dcache_io_ptw_pmp_6_addr; // @[HellaCache.scala 215:43]
  wire [31:0] dcache_io_ptw_pmp_6_mask; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_7_cfg_l; // @[HellaCache.scala 215:43]
  wire [1:0] dcache_io_ptw_pmp_7_cfg_a; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_7_cfg_x; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_7_cfg_w; // @[HellaCache.scala 215:43]
  wire  dcache_io_ptw_pmp_7_cfg_r; // @[HellaCache.scala 215:43]
  wire [29:0] dcache_io_ptw_pmp_7_addr; // @[HellaCache.scala 215:43]
  wire [31:0] dcache_io_ptw_pmp_7_mask; // @[HellaCache.scala 215:43]
  wire [26:0] dcache_io_ptw_vpoffset_bits_value; // @[HellaCache.scala 215:43]
  wire [29:0] dcache_io_covSum; // @[HellaCache.scala 215:43]
  wire  dcache_metaAssert; // @[HellaCache.scala 215:43]
  wire  dcache_metaReset; // @[HellaCache.scala 215:43]
  wire  dcache_data_halt; // @[HellaCache.scala 215:43]
  wire  dcache_tlb_halt; // @[HellaCache.scala 215:43]
  wire  frontend_gated_clock; // @[Frontend.scala 340:28]
  wire  frontend_reset; // @[Frontend.scala 340:28]
  wire  frontend_auto_icache_master_out_a_ready; // @[Frontend.scala 340:28]
  wire  frontend_auto_icache_master_out_a_valid; // @[Frontend.scala 340:28]
  wire [31:0] frontend_auto_icache_master_out_a_bits_address; // @[Frontend.scala 340:28]
  wire  frontend_auto_icache_master_out_d_valid; // @[Frontend.scala 340:28]
  wire [2:0] frontend_auto_icache_master_out_d_bits_opcode; // @[Frontend.scala 340:28]
  wire [3:0] frontend_auto_icache_master_out_d_bits_size; // @[Frontend.scala 340:28]
  wire [63:0] frontend_auto_icache_master_out_d_bits_data; // @[Frontend.scala 340:28]
  wire  frontend_auto_icache_master_out_d_bits_corrupt; // @[Frontend.scala 340:28]
  wire [31:0] frontend_io_reset_vector; // @[Frontend.scala 340:28]
  wire  frontend_io_cpu_might_request; // @[Frontend.scala 340:28]
  wire  frontend_io_cpu_req_valid; // @[Frontend.scala 340:28]
  wire [39:0] frontend_io_cpu_req_bits_pc; // @[Frontend.scala 340:28]
  wire  frontend_io_cpu_req_bits_speculative; // @[Frontend.scala 340:28]
  wire  frontend_io_cpu_sfence_valid; // @[Frontend.scala 340:28]
  wire  frontend_io_cpu_sfence_bits_rs1; // @[Frontend.scala 340:28]
  wire  frontend_io_cpu_sfence_bits_rs2; // @[Frontend.scala 340:28]
  wire [38:0] frontend_io_cpu_sfence_bits_addr; // @[Frontend.scala 340:28]
  wire  frontend_io_cpu_resp_ready; // @[Frontend.scala 340:28]
  wire  frontend_io_cpu_resp_valid; // @[Frontend.scala 340:28]
  wire  frontend_io_cpu_resp_bits_btb_taken; // @[Frontend.scala 340:28]
  wire  frontend_io_cpu_resp_bits_btb_bridx; // @[Frontend.scala 340:28]
  wire [4:0] frontend_io_cpu_resp_bits_btb_entry; // @[Frontend.scala 340:28]
  wire [7:0] frontend_io_cpu_resp_bits_btb_bht_history; // @[Frontend.scala 340:28]
  wire [39:0] frontend_io_cpu_resp_bits_pc; // @[Frontend.scala 340:28]
  wire [31:0] frontend_io_cpu_resp_bits_data; // @[Frontend.scala 340:28]
  wire  frontend_io_cpu_resp_bits_xcpt_pf_inst; // @[Frontend.scala 340:28]
  wire  frontend_io_cpu_resp_bits_xcpt_ae_inst; // @[Frontend.scala 340:28]
  wire  frontend_io_cpu_resp_bits_replay; // @[Frontend.scala 340:28]
  wire  frontend_io_cpu_btb_update_valid; // @[Frontend.scala 340:28]
  wire [4:0] frontend_io_cpu_btb_update_bits_prediction_entry; // @[Frontend.scala 340:28]
  wire [38:0] frontend_io_cpu_btb_update_bits_pc; // @[Frontend.scala 340:28]
  wire  frontend_io_cpu_btb_update_bits_isValid; // @[Frontend.scala 340:28]
  wire [38:0] frontend_io_cpu_btb_update_bits_br_pc; // @[Frontend.scala 340:28]
  wire [1:0] frontend_io_cpu_btb_update_bits_cfiType; // @[Frontend.scala 340:28]
  wire  frontend_io_cpu_bht_update_valid; // @[Frontend.scala 340:28]
  wire [7:0] frontend_io_cpu_bht_update_bits_prediction_history; // @[Frontend.scala 340:28]
  wire [38:0] frontend_io_cpu_bht_update_bits_pc; // @[Frontend.scala 340:28]
  wire  frontend_io_cpu_bht_update_bits_branch; // @[Frontend.scala 340:28]
  wire  frontend_io_cpu_bht_update_bits_taken; // @[Frontend.scala 340:28]
  wire  frontend_io_cpu_bht_update_bits_mispredict; // @[Frontend.scala 340:28]
  wire  frontend_io_cpu_flush_icache; // @[Frontend.scala 340:28]
  wire [39:0] frontend_io_cpu_npc; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_req_ready; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_req_valid; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_req_bits_valid; // @[Frontend.scala 340:28]
  wire [26:0] frontend_io_ptw_req_bits_bits_addr; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_resp_valid; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_resp_bits_ae; // @[Frontend.scala 340:28]
  wire [53:0] frontend_io_ptw_resp_bits_pte_ppn; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_resp_bits_pte_d; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_resp_bits_pte_a; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_resp_bits_pte_g; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_resp_bits_pte_u; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_resp_bits_pte_x; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_resp_bits_pte_w; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_resp_bits_pte_r; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_resp_bits_pte_v; // @[Frontend.scala 340:28]
  wire [1:0] frontend_io_ptw_resp_bits_level; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_resp_bits_homogeneous; // @[Frontend.scala 340:28]
  wire [3:0] frontend_io_ptw_ptbr_mode; // @[Frontend.scala 340:28]
  wire [1:0] frontend_io_ptw_status_prv; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_0_cfg_l; // @[Frontend.scala 340:28]
  wire [1:0] frontend_io_ptw_pmp_0_cfg_a; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_0_cfg_x; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_0_cfg_w; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_0_cfg_r; // @[Frontend.scala 340:28]
  wire [29:0] frontend_io_ptw_pmp_0_addr; // @[Frontend.scala 340:28]
  wire [31:0] frontend_io_ptw_pmp_0_mask; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_1_cfg_l; // @[Frontend.scala 340:28]
  wire [1:0] frontend_io_ptw_pmp_1_cfg_a; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_1_cfg_x; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_1_cfg_w; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_1_cfg_r; // @[Frontend.scala 340:28]
  wire [29:0] frontend_io_ptw_pmp_1_addr; // @[Frontend.scala 340:28]
  wire [31:0] frontend_io_ptw_pmp_1_mask; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_2_cfg_l; // @[Frontend.scala 340:28]
  wire [1:0] frontend_io_ptw_pmp_2_cfg_a; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_2_cfg_x; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_2_cfg_w; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_2_cfg_r; // @[Frontend.scala 340:28]
  wire [29:0] frontend_io_ptw_pmp_2_addr; // @[Frontend.scala 340:28]
  wire [31:0] frontend_io_ptw_pmp_2_mask; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_3_cfg_l; // @[Frontend.scala 340:28]
  wire [1:0] frontend_io_ptw_pmp_3_cfg_a; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_3_cfg_x; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_3_cfg_w; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_3_cfg_r; // @[Frontend.scala 340:28]
  wire [29:0] frontend_io_ptw_pmp_3_addr; // @[Frontend.scala 340:28]
  wire [31:0] frontend_io_ptw_pmp_3_mask; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_4_cfg_l; // @[Frontend.scala 340:28]
  wire [1:0] frontend_io_ptw_pmp_4_cfg_a; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_4_cfg_x; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_4_cfg_w; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_4_cfg_r; // @[Frontend.scala 340:28]
  wire [29:0] frontend_io_ptw_pmp_4_addr; // @[Frontend.scala 340:28]
  wire [31:0] frontend_io_ptw_pmp_4_mask; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_5_cfg_l; // @[Frontend.scala 340:28]
  wire [1:0] frontend_io_ptw_pmp_5_cfg_a; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_5_cfg_x; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_5_cfg_w; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_5_cfg_r; // @[Frontend.scala 340:28]
  wire [29:0] frontend_io_ptw_pmp_5_addr; // @[Frontend.scala 340:28]
  wire [31:0] frontend_io_ptw_pmp_5_mask; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_6_cfg_l; // @[Frontend.scala 340:28]
  wire [1:0] frontend_io_ptw_pmp_6_cfg_a; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_6_cfg_x; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_6_cfg_w; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_6_cfg_r; // @[Frontend.scala 340:28]
  wire [29:0] frontend_io_ptw_pmp_6_addr; // @[Frontend.scala 340:28]
  wire [31:0] frontend_io_ptw_pmp_6_mask; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_7_cfg_l; // @[Frontend.scala 340:28]
  wire [1:0] frontend_io_ptw_pmp_7_cfg_a; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_7_cfg_x; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_7_cfg_w; // @[Frontend.scala 340:28]
  wire  frontend_io_ptw_pmp_7_cfg_r; // @[Frontend.scala 340:28]
  wire [29:0] frontend_io_ptw_pmp_7_addr; // @[Frontend.scala 340:28]
  wire [31:0] frontend_io_ptw_pmp_7_mask; // @[Frontend.scala 340:28]
  wire [26:0] frontend_io_ptw_vpoffset_bits_value; // @[Frontend.scala 340:28]
  wire [29:0] frontend_io_covSum; // @[Frontend.scala 340:28]
  wire  frontend_metaAssert; // @[Frontend.scala 340:28]
  wire  frontend_metaReset; // @[Frontend.scala 340:28]
  wire  frontend_icache_halt; // @[Frontend.scala 340:28]
  wire  frontend_fq_halt; // @[Frontend.scala 340:28]
  wire  frontend_tlb_halt; // @[Frontend.scala 340:28]
  wire  frontend_btb_halt; // @[Frontend.scala 340:28]
  wire  buffer_clock; // @[Buffer.scala 69:28]
  wire  buffer_reset; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_a_ready; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_a_valid; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_a_bits_opcode; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_a_bits_param; // @[Buffer.scala 69:28]
  wire [3:0] buffer_auto_in_a_bits_size; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_a_bits_source; // @[Buffer.scala 69:28]
  wire [31:0] buffer_auto_in_a_bits_address; // @[Buffer.scala 69:28]
  wire [7:0] buffer_auto_in_a_bits_mask; // @[Buffer.scala 69:28]
  wire [63:0] buffer_auto_in_a_bits_data; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_a_bits_corrupt; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_b_ready; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_b_valid; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_b_bits_opcode; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_b_bits_param; // @[Buffer.scala 69:28]
  wire [3:0] buffer_auto_in_b_bits_size; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_b_bits_source; // @[Buffer.scala 69:28]
  wire [31:0] buffer_auto_in_b_bits_address; // @[Buffer.scala 69:28]
  wire [7:0] buffer_auto_in_b_bits_mask; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_b_bits_corrupt; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_c_ready; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_c_valid; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_c_bits_opcode; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_c_bits_param; // @[Buffer.scala 69:28]
  wire [3:0] buffer_auto_in_c_bits_size; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_c_bits_source; // @[Buffer.scala 69:28]
  wire [31:0] buffer_auto_in_c_bits_address; // @[Buffer.scala 69:28]
  wire [63:0] buffer_auto_in_c_bits_data; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_d_ready; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_d_valid; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_d_bits_opcode; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_d_bits_param; // @[Buffer.scala 69:28]
  wire [3:0] buffer_auto_in_d_bits_size; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_d_bits_source; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_d_bits_sink; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_d_bits_denied; // @[Buffer.scala 69:28]
  wire [63:0] buffer_auto_in_d_bits_data; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_d_bits_corrupt; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_e_ready; // @[Buffer.scala 69:28]
  wire  buffer_auto_in_e_valid; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_e_bits_sink; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_a_ready; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_a_valid; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_a_bits_opcode; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_a_bits_param; // @[Buffer.scala 69:28]
  wire [3:0] buffer_auto_out_a_bits_size; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_a_bits_source; // @[Buffer.scala 69:28]
  wire [31:0] buffer_auto_out_a_bits_address; // @[Buffer.scala 69:28]
  wire [7:0] buffer_auto_out_a_bits_mask; // @[Buffer.scala 69:28]
  wire [63:0] buffer_auto_out_a_bits_data; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_a_bits_corrupt; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_b_ready; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_b_valid; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_b_bits_opcode; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_b_bits_param; // @[Buffer.scala 69:28]
  wire [3:0] buffer_auto_out_b_bits_size; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_b_bits_source; // @[Buffer.scala 69:28]
  wire [31:0] buffer_auto_out_b_bits_address; // @[Buffer.scala 69:28]
  wire [7:0] buffer_auto_out_b_bits_mask; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_b_bits_corrupt; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_c_ready; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_c_valid; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_c_bits_opcode; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_c_bits_param; // @[Buffer.scala 69:28]
  wire [3:0] buffer_auto_out_c_bits_size; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_c_bits_source; // @[Buffer.scala 69:28]
  wire [31:0] buffer_auto_out_c_bits_address; // @[Buffer.scala 69:28]
  wire [63:0] buffer_auto_out_c_bits_data; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_c_bits_corrupt; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_d_ready; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_d_valid; // @[Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_d_bits_opcode; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_d_bits_param; // @[Buffer.scala 69:28]
  wire [3:0] buffer_auto_out_d_bits_size; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_d_bits_source; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_d_bits_sink; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_d_bits_denied; // @[Buffer.scala 69:28]
  wire [63:0] buffer_auto_out_d_bits_data; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_d_bits_corrupt; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_e_ready; // @[Buffer.scala 69:28]
  wire  buffer_auto_out_e_valid; // @[Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_e_bits_sink; // @[Buffer.scala 69:28]
  wire [29:0] buffer_io_covSum; // @[Buffer.scala 69:28]
  wire  buffer_metaAssert; // @[Buffer.scala 69:28]
  wire  buffer_metaReset; // @[Buffer.scala 69:28]
  wire  buffer_TLMonitor_halt; // @[Buffer.scala 69:28]
  wire  buffer_Queue_4_halt; // @[Buffer.scala 69:28]
  wire  buffer_Queue_2_halt; // @[Buffer.scala 69:28]
  wire  buffer_Queue_1_halt; // @[Buffer.scala 69:28]
  wire  buffer_Queue_3_halt; // @[Buffer.scala 69:28]
  wire  buffer_Queue_halt; // @[Buffer.scala 69:28]
  wire  intsink_clock; // @[Crossing.scala 63:29]
  wire  intsink_auto_in_sync_0; // @[Crossing.scala 63:29]
  wire  intsink_auto_out_0; // @[Crossing.scala 63:29]
  wire [29:0] intsink_io_covSum; // @[Crossing.scala 63:29]
  wire  intsink_metaAssert; // @[Crossing.scala 63:29]
  wire  intsink_metaReset; // @[Crossing.scala 63:29]
  wire  intsink_SynchronizerShiftReg_w1_d3_halt; // @[Crossing.scala 63:29]
  wire  intsink_1_auto_in_sync_0; // @[Crossing.scala 63:29]
  wire  intsink_1_auto_in_sync_1; // @[Crossing.scala 63:29]
  wire  intsink_1_auto_out_0; // @[Crossing.scala 63:29]
  wire  intsink_1_auto_out_1; // @[Crossing.scala 63:29]
  wire [29:0] intsink_1_io_covSum; // @[Crossing.scala 63:29]
  wire  intsink_1_metaAssert; // @[Crossing.scala 63:29]
  wire  intsink_2_auto_in_sync_0; // @[Crossing.scala 63:29]
  wire  intsink_2_auto_out_0; // @[Crossing.scala 63:29]
  wire [29:0] intsink_2_io_covSum; // @[Crossing.scala 63:29]
  wire  intsink_2_metaAssert; // @[Crossing.scala 63:29]
  wire  intsink_3_auto_in_sync_0; // @[Crossing.scala 63:29]
  wire  intsink_3_auto_out_0; // @[Crossing.scala 63:29]
  wire [29:0] intsink_3_io_covSum; // @[Crossing.scala 63:29]
  wire  intsink_3_metaAssert; // @[Crossing.scala 63:29]
  wire  fpuOpt_clock; // @[RocketTile.scala 173:62]
  wire  fpuOpt_reset; // @[RocketTile.scala 173:62]
  wire [31:0] fpuOpt_io_inst; // @[RocketTile.scala 173:62]
  wire [63:0] fpuOpt_io_fromint_data; // @[RocketTile.scala 173:62]
  wire [2:0] fpuOpt_io_fcsr_rm; // @[RocketTile.scala 173:62]
  wire  fpuOpt_io_fcsr_flags_valid; // @[RocketTile.scala 173:62]
  wire [4:0] fpuOpt_io_fcsr_flags_bits; // @[RocketTile.scala 173:62]
  wire [63:0] fpuOpt_io_store_data; // @[RocketTile.scala 173:62]
  wire [63:0] fpuOpt_io_toint_data; // @[RocketTile.scala 173:62]
  wire  fpuOpt_io_dmem_resp_val; // @[RocketTile.scala 173:62]
  wire [2:0] fpuOpt_io_dmem_resp_type; // @[RocketTile.scala 173:62]
  wire [4:0] fpuOpt_io_dmem_resp_tag; // @[RocketTile.scala 173:62]
  wire [63:0] fpuOpt_io_dmem_resp_data; // @[RocketTile.scala 173:62]
  wire  fpuOpt_io_valid; // @[RocketTile.scala 173:62]
  wire  fpuOpt_io_fcsr_rdy; // @[RocketTile.scala 173:62]
  wire  fpuOpt_io_nack_mem; // @[RocketTile.scala 173:62]
  wire  fpuOpt_io_illegal_rm; // @[RocketTile.scala 173:62]
  wire  fpuOpt_io_killx; // @[RocketTile.scala 173:62]
  wire  fpuOpt_io_killm; // @[RocketTile.scala 173:62]
  wire  fpuOpt_io_dec_wen; // @[RocketTile.scala 173:62]
  wire  fpuOpt_io_dec_ren1; // @[RocketTile.scala 173:62]
  wire  fpuOpt_io_dec_ren2; // @[RocketTile.scala 173:62]
  wire  fpuOpt_io_dec_ren3; // @[RocketTile.scala 173:62]
  wire  fpuOpt_io_sboard_set; // @[RocketTile.scala 173:62]
  wire  fpuOpt_io_sboard_clr; // @[RocketTile.scala 173:62]
  wire [4:0] fpuOpt_io_sboard_clra; // @[RocketTile.scala 173:62]
  wire [29:0] fpuOpt_io_covSum; // @[RocketTile.scala 173:62]
  wire  fpuOpt_metaAssert; // @[RocketTile.scala 173:62]
  wire  fpuOpt_metaReset; // @[RocketTile.scala 173:62]
  wire  fpuOpt_dfma_halt; // @[RocketTile.scala 173:62]
  wire  fpuOpt_fpmu_halt; // @[RocketTile.scala 173:62]
  wire  fpuOpt_divSqrt_1_halt; // @[RocketTile.scala 173:62]
  wire  fpuOpt_ifpu_halt; // @[RocketTile.scala 173:62]
  wire  fpuOpt_divSqrt_halt; // @[RocketTile.scala 173:62]
  wire  fpuOpt_fpiu_halt; // @[RocketTile.scala 173:62]
  wire  fpuOpt_sfma_halt; // @[RocketTile.scala 173:62]
  wire  dcacheArb_clock; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_0_req_ready; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_0_req_valid; // @[HellaCache.scala 227:25]
  wire [39:0] dcacheArb_io_requestor_0_req_bits_addr; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_0_s1_kill; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_0_s2_nack; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_0_resp_valid; // @[HellaCache.scala 227:25]
  wire [63:0] dcacheArb_io_requestor_0_resp_bits_data_word_bypass; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_0_s2_xcpt_ae_ld; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_1_req_ready; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_1_req_valid; // @[HellaCache.scala 227:25]
  wire [39:0] dcacheArb_io_requestor_1_req_bits_addr; // @[HellaCache.scala 227:25]
  wire [6:0] dcacheArb_io_requestor_1_req_bits_tag; // @[HellaCache.scala 227:25]
  wire [4:0] dcacheArb_io_requestor_1_req_bits_cmd; // @[HellaCache.scala 227:25]
  wire [2:0] dcacheArb_io_requestor_1_req_bits_typ; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_1_s1_kill; // @[HellaCache.scala 227:25]
  wire [63:0] dcacheArb_io_requestor_1_s1_data_data; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_1_s2_nack; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_1_resp_valid; // @[HellaCache.scala 227:25]
  wire [6:0] dcacheArb_io_requestor_1_resp_bits_tag; // @[HellaCache.scala 227:25]
  wire [2:0] dcacheArb_io_requestor_1_resp_bits_typ; // @[HellaCache.scala 227:25]
  wire [63:0] dcacheArb_io_requestor_1_resp_bits_data; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_1_resp_bits_replay; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_1_resp_bits_has_data; // @[HellaCache.scala 227:25]
  wire [63:0] dcacheArb_io_requestor_1_resp_bits_data_word_bypass; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_1_replay_next; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_ma_ld; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_ma_st; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_pf_ld; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_pf_st; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_ae_ld; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_ae_st; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_1_ordered; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_1_perf_grant; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_1_keep_clock_enabled; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_requestor_1_clock_enabled; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_mem_req_ready; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_mem_req_valid; // @[HellaCache.scala 227:25]
  wire [39:0] dcacheArb_io_mem_req_bits_addr; // @[HellaCache.scala 227:25]
  wire [6:0] dcacheArb_io_mem_req_bits_tag; // @[HellaCache.scala 227:25]
  wire [4:0] dcacheArb_io_mem_req_bits_cmd; // @[HellaCache.scala 227:25]
  wire [2:0] dcacheArb_io_mem_req_bits_typ; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_mem_req_bits_phys; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_mem_s1_kill; // @[HellaCache.scala 227:25]
  wire [63:0] dcacheArb_io_mem_s1_data_data; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_mem_s2_nack; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_mem_resp_valid; // @[HellaCache.scala 227:25]
  wire [6:0] dcacheArb_io_mem_resp_bits_tag; // @[HellaCache.scala 227:25]
  wire [2:0] dcacheArb_io_mem_resp_bits_typ; // @[HellaCache.scala 227:25]
  wire [63:0] dcacheArb_io_mem_resp_bits_data; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_mem_resp_bits_replay; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_mem_resp_bits_has_data; // @[HellaCache.scala 227:25]
  wire [63:0] dcacheArb_io_mem_resp_bits_data_word_bypass; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_mem_replay_next; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_mem_s2_xcpt_ma_ld; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_mem_s2_xcpt_ma_st; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_mem_s2_xcpt_pf_ld; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_mem_s2_xcpt_pf_st; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_mem_s2_xcpt_ae_ld; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_mem_s2_xcpt_ae_st; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_mem_ordered; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_mem_perf_grant; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_mem_keep_clock_enabled; // @[HellaCache.scala 227:25]
  wire  dcacheArb_io_mem_clock_enabled; // @[HellaCache.scala 227:25]
  wire [29:0] dcacheArb_io_covSum; // @[HellaCache.scala 227:25]
  wire  dcacheArb_metaAssert; // @[HellaCache.scala 227:25]
  wire  dcacheArb_metaReset; // @[HellaCache.scala 227:25]
  wire  ptw_clock; // @[PTW.scala 531:19]
  wire  ptw_reset; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_req_ready; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_req_valid; // @[PTW.scala 531:19]
  wire [26:0] ptw_io_requestor_0_req_bits_bits_addr; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_resp_valid; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_resp_bits_ae; // @[PTW.scala 531:19]
  wire [53:0] ptw_io_requestor_0_resp_bits_pte_ppn; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_resp_bits_pte_d; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_resp_bits_pte_a; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_resp_bits_pte_g; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_resp_bits_pte_u; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_resp_bits_pte_x; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_resp_bits_pte_w; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_resp_bits_pte_r; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_resp_bits_pte_v; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_requestor_0_resp_bits_level; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_resp_bits_homogeneous; // @[PTW.scala 531:19]
  wire [3:0] ptw_io_requestor_0_ptbr_mode; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_requestor_0_status_dprv; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_status_mxr; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_status_sum; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_0_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_requestor_0_pmp_0_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_0_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_0_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_0_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_requestor_0_pmp_0_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_requestor_0_pmp_0_mask; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_1_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_requestor_0_pmp_1_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_1_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_1_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_1_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_requestor_0_pmp_1_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_requestor_0_pmp_1_mask; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_2_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_requestor_0_pmp_2_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_2_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_2_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_2_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_requestor_0_pmp_2_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_requestor_0_pmp_2_mask; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_3_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_requestor_0_pmp_3_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_3_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_3_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_3_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_requestor_0_pmp_3_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_requestor_0_pmp_3_mask; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_4_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_requestor_0_pmp_4_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_4_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_4_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_4_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_requestor_0_pmp_4_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_requestor_0_pmp_4_mask; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_5_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_requestor_0_pmp_5_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_5_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_5_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_5_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_requestor_0_pmp_5_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_requestor_0_pmp_5_mask; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_6_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_requestor_0_pmp_6_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_6_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_6_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_6_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_requestor_0_pmp_6_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_requestor_0_pmp_6_mask; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_7_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_requestor_0_pmp_7_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_7_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_7_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_0_pmp_7_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_requestor_0_pmp_7_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_requestor_0_pmp_7_mask; // @[PTW.scala 531:19]
  wire [26:0] ptw_io_requestor_0_vpoffset_bits_value; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_req_ready; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_req_valid; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_req_bits_valid; // @[PTW.scala 531:19]
  wire [26:0] ptw_io_requestor_1_req_bits_bits_addr; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_resp_valid; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_resp_bits_ae; // @[PTW.scala 531:19]
  wire [53:0] ptw_io_requestor_1_resp_bits_pte_ppn; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_resp_bits_pte_d; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_resp_bits_pte_a; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_resp_bits_pte_g; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_resp_bits_pte_u; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_resp_bits_pte_x; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_resp_bits_pte_w; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_resp_bits_pte_r; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_resp_bits_pte_v; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_requestor_1_resp_bits_level; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_resp_bits_homogeneous; // @[PTW.scala 531:19]
  wire [3:0] ptw_io_requestor_1_ptbr_mode; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_requestor_1_status_prv; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_0_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_requestor_1_pmp_0_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_0_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_0_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_0_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_requestor_1_pmp_0_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_requestor_1_pmp_0_mask; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_1_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_requestor_1_pmp_1_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_1_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_1_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_1_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_requestor_1_pmp_1_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_requestor_1_pmp_1_mask; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_2_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_requestor_1_pmp_2_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_2_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_2_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_2_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_requestor_1_pmp_2_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_requestor_1_pmp_2_mask; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_3_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_requestor_1_pmp_3_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_3_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_3_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_3_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_requestor_1_pmp_3_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_requestor_1_pmp_3_mask; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_4_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_requestor_1_pmp_4_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_4_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_4_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_4_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_requestor_1_pmp_4_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_requestor_1_pmp_4_mask; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_5_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_requestor_1_pmp_5_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_5_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_5_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_5_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_requestor_1_pmp_5_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_requestor_1_pmp_5_mask; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_6_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_requestor_1_pmp_6_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_6_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_6_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_6_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_requestor_1_pmp_6_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_requestor_1_pmp_6_mask; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_7_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_requestor_1_pmp_7_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_7_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_7_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_requestor_1_pmp_7_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_requestor_1_pmp_7_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_requestor_1_pmp_7_mask; // @[PTW.scala 531:19]
  wire [26:0] ptw_io_requestor_1_vpoffset_bits_value; // @[PTW.scala 531:19]
  wire  ptw_io_mem_req_ready; // @[PTW.scala 531:19]
  wire  ptw_io_mem_req_valid; // @[PTW.scala 531:19]
  wire [39:0] ptw_io_mem_req_bits_addr; // @[PTW.scala 531:19]
  wire  ptw_io_mem_s1_kill; // @[PTW.scala 531:19]
  wire  ptw_io_mem_s2_nack; // @[PTW.scala 531:19]
  wire  ptw_io_mem_resp_valid; // @[PTW.scala 531:19]
  wire [63:0] ptw_io_mem_resp_bits_data_word_bypass; // @[PTW.scala 531:19]
  wire  ptw_io_mem_s2_xcpt_ae_ld; // @[PTW.scala 531:19]
  wire [3:0] ptw_io_dpath_ptbr_mode; // @[PTW.scala 531:19]
  wire [43:0] ptw_io_dpath_ptbr_ppn; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_sfence_valid; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_sfence_bits_rs1; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_dpath_status_dprv; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_dpath_status_prv; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_status_mxr; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_status_sum; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_0_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_dpath_pmp_0_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_0_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_0_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_0_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_dpath_pmp_0_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_dpath_pmp_0_mask; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_1_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_dpath_pmp_1_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_1_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_1_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_1_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_dpath_pmp_1_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_dpath_pmp_1_mask; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_2_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_dpath_pmp_2_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_2_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_2_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_2_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_dpath_pmp_2_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_dpath_pmp_2_mask; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_3_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_dpath_pmp_3_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_3_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_3_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_3_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_dpath_pmp_3_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_dpath_pmp_3_mask; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_4_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_dpath_pmp_4_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_4_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_4_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_4_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_dpath_pmp_4_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_dpath_pmp_4_mask; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_5_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_dpath_pmp_5_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_5_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_5_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_5_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_dpath_pmp_5_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_dpath_pmp_5_mask; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_6_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_dpath_pmp_6_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_6_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_6_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_6_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_dpath_pmp_6_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_dpath_pmp_6_mask; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_7_cfg_l; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_dpath_pmp_7_cfg_a; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_7_cfg_x; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_7_cfg_w; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pmp_7_cfg_r; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_dpath_pmp_7_addr; // @[PTW.scala 531:19]
  wire [31:0] ptw_io_dpath_pmp_7_mask; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pcode_req_valid; // @[PTW.scala 531:19]
  wire [1:0] ptw_io_dpath_pcode_req_bits_id; // @[PTW.scala 531:19]
  wire [19:0] ptw_io_dpath_pcode_req_bits_value_base; // @[PTW.scala 531:19]
  wire [9:0] ptw_io_dpath_pcode_req_bits_value_mask; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pcode_req_bits_value_valid; // @[PTW.scala 531:19]
  wire  ptw_io_dpath_pcode_req_bits_value_locked; // @[PTW.scala 531:19]
  wire [26:0] ptw_io_dpath_vpoffset_req_bits_value; // @[PTW.scala 531:19]
  wire [29:0] ptw_io_covSum; // @[PTW.scala 531:19]
  wire  ptw_metaAssert; // @[PTW.scala 531:19]
  wire  ptw_metaReset; // @[PTW.scala 531:19]
  wire  ptw_arb_halt; // @[PTW.scala 531:19]
  wire  core_clock; // @[RocketTile.scala 115:20]
  wire  core_reset; // @[RocketTile.scala 115:20]
  wire [1:0] core_io_hartid; // @[RocketTile.scala 115:20]
  wire  core_io_interrupts_debug; // @[RocketTile.scala 115:20]
  wire  core_io_interrupts_mtip; // @[RocketTile.scala 115:20]
  wire  core_io_interrupts_msip; // @[RocketTile.scala 115:20]
  wire  core_io_interrupts_meip; // @[RocketTile.scala 115:20]
  wire  core_io_interrupts_seip; // @[RocketTile.scala 115:20]
  wire  core_io_imem_might_request; // @[RocketTile.scala 115:20]
  wire  core_io_imem_req_valid; // @[RocketTile.scala 115:20]
  wire [39:0] core_io_imem_req_bits_pc; // @[RocketTile.scala 115:20]
  wire  core_io_imem_req_bits_speculative; // @[RocketTile.scala 115:20]
  wire  core_io_imem_sfence_valid; // @[RocketTile.scala 115:20]
  wire  core_io_imem_sfence_bits_rs1; // @[RocketTile.scala 115:20]
  wire  core_io_imem_sfence_bits_rs2; // @[RocketTile.scala 115:20]
  wire [38:0] core_io_imem_sfence_bits_addr; // @[RocketTile.scala 115:20]
  wire  core_io_imem_resp_ready; // @[RocketTile.scala 115:20]
  wire  core_io_imem_resp_valid; // @[RocketTile.scala 115:20]
  wire  core_io_imem_resp_bits_btb_taken; // @[RocketTile.scala 115:20]
  wire  core_io_imem_resp_bits_btb_bridx; // @[RocketTile.scala 115:20]
  wire [4:0] core_io_imem_resp_bits_btb_entry; // @[RocketTile.scala 115:20]
  wire [7:0] core_io_imem_resp_bits_btb_bht_history; // @[RocketTile.scala 115:20]
  wire [39:0] core_io_imem_resp_bits_pc; // @[RocketTile.scala 115:20]
  wire [31:0] core_io_imem_resp_bits_data; // @[RocketTile.scala 115:20]
  wire  core_io_imem_resp_bits_xcpt_pf_inst; // @[RocketTile.scala 115:20]
  wire  core_io_imem_resp_bits_xcpt_ae_inst; // @[RocketTile.scala 115:20]
  wire  core_io_imem_resp_bits_replay; // @[RocketTile.scala 115:20]
  wire  core_io_imem_btb_update_valid; // @[RocketTile.scala 115:20]
  wire [4:0] core_io_imem_btb_update_bits_prediction_entry; // @[RocketTile.scala 115:20]
  wire [38:0] core_io_imem_btb_update_bits_pc; // @[RocketTile.scala 115:20]
  wire  core_io_imem_btb_update_bits_isValid; // @[RocketTile.scala 115:20]
  wire [38:0] core_io_imem_btb_update_bits_br_pc; // @[RocketTile.scala 115:20]
  wire [1:0] core_io_imem_btb_update_bits_cfiType; // @[RocketTile.scala 115:20]
  wire  core_io_imem_bht_update_valid; // @[RocketTile.scala 115:20]
  wire [7:0] core_io_imem_bht_update_bits_prediction_history; // @[RocketTile.scala 115:20]
  wire [38:0] core_io_imem_bht_update_bits_pc; // @[RocketTile.scala 115:20]
  wire  core_io_imem_bht_update_bits_branch; // @[RocketTile.scala 115:20]
  wire  core_io_imem_bht_update_bits_taken; // @[RocketTile.scala 115:20]
  wire  core_io_imem_bht_update_bits_mispredict; // @[RocketTile.scala 115:20]
  wire  core_io_imem_flush_icache; // @[RocketTile.scala 115:20]
  wire  core_io_dmem_req_ready; // @[RocketTile.scala 115:20]
  wire  core_io_dmem_req_valid; // @[RocketTile.scala 115:20]
  wire [39:0] core_io_dmem_req_bits_addr; // @[RocketTile.scala 115:20]
  wire [6:0] core_io_dmem_req_bits_tag; // @[RocketTile.scala 115:20]
  wire [4:0] core_io_dmem_req_bits_cmd; // @[RocketTile.scala 115:20]
  wire [2:0] core_io_dmem_req_bits_typ; // @[RocketTile.scala 115:20]
  wire  core_io_dmem_s1_kill; // @[RocketTile.scala 115:20]
  wire [63:0] core_io_dmem_s1_data_data; // @[RocketTile.scala 115:20]
  wire  core_io_dmem_s2_nack; // @[RocketTile.scala 115:20]
  wire  core_io_dmem_resp_valid; // @[RocketTile.scala 115:20]
  wire [6:0] core_io_dmem_resp_bits_tag; // @[RocketTile.scala 115:20]
  wire [2:0] core_io_dmem_resp_bits_typ; // @[RocketTile.scala 115:20]
  wire [63:0] core_io_dmem_resp_bits_data; // @[RocketTile.scala 115:20]
  wire  core_io_dmem_resp_bits_replay; // @[RocketTile.scala 115:20]
  wire  core_io_dmem_resp_bits_has_data; // @[RocketTile.scala 115:20]
  wire [63:0] core_io_dmem_resp_bits_data_word_bypass; // @[RocketTile.scala 115:20]
  wire  core_io_dmem_replay_next; // @[RocketTile.scala 115:20]
  wire  core_io_dmem_s2_xcpt_ma_ld; // @[RocketTile.scala 115:20]
  wire  core_io_dmem_s2_xcpt_ma_st; // @[RocketTile.scala 115:20]
  wire  core_io_dmem_s2_xcpt_pf_ld; // @[RocketTile.scala 115:20]
  wire  core_io_dmem_s2_xcpt_pf_st; // @[RocketTile.scala 115:20]
  wire  core_io_dmem_s2_xcpt_ae_ld; // @[RocketTile.scala 115:20]
  wire  core_io_dmem_s2_xcpt_ae_st; // @[RocketTile.scala 115:20]
  wire  core_io_dmem_ordered; // @[RocketTile.scala 115:20]
  wire  core_io_dmem_perf_grant; // @[RocketTile.scala 115:20]
  wire  core_io_dmem_keep_clock_enabled; // @[RocketTile.scala 115:20]
  wire  core_io_dmem_clock_enabled; // @[RocketTile.scala 115:20]
  wire [3:0] core_io_ptw_ptbr_mode; // @[RocketTile.scala 115:20]
  wire [43:0] core_io_ptw_ptbr_ppn; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_sfence_valid; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_sfence_bits_rs1; // @[RocketTile.scala 115:20]
  wire [1:0] core_io_ptw_status_dprv; // @[RocketTile.scala 115:20]
  wire [1:0] core_io_ptw_status_prv; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_status_mxr; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_status_sum; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_0_cfg_l; // @[RocketTile.scala 115:20]
  wire [1:0] core_io_ptw_pmp_0_cfg_a; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_0_cfg_x; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_0_cfg_w; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_0_cfg_r; // @[RocketTile.scala 115:20]
  wire [29:0] core_io_ptw_pmp_0_addr; // @[RocketTile.scala 115:20]
  wire [31:0] core_io_ptw_pmp_0_mask; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_1_cfg_l; // @[RocketTile.scala 115:20]
  wire [1:0] core_io_ptw_pmp_1_cfg_a; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_1_cfg_x; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_1_cfg_w; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_1_cfg_r; // @[RocketTile.scala 115:20]
  wire [29:0] core_io_ptw_pmp_1_addr; // @[RocketTile.scala 115:20]
  wire [31:0] core_io_ptw_pmp_1_mask; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_2_cfg_l; // @[RocketTile.scala 115:20]
  wire [1:0] core_io_ptw_pmp_2_cfg_a; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_2_cfg_x; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_2_cfg_w; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_2_cfg_r; // @[RocketTile.scala 115:20]
  wire [29:0] core_io_ptw_pmp_2_addr; // @[RocketTile.scala 115:20]
  wire [31:0] core_io_ptw_pmp_2_mask; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_3_cfg_l; // @[RocketTile.scala 115:20]
  wire [1:0] core_io_ptw_pmp_3_cfg_a; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_3_cfg_x; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_3_cfg_w; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_3_cfg_r; // @[RocketTile.scala 115:20]
  wire [29:0] core_io_ptw_pmp_3_addr; // @[RocketTile.scala 115:20]
  wire [31:0] core_io_ptw_pmp_3_mask; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_4_cfg_l; // @[RocketTile.scala 115:20]
  wire [1:0] core_io_ptw_pmp_4_cfg_a; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_4_cfg_x; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_4_cfg_w; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_4_cfg_r; // @[RocketTile.scala 115:20]
  wire [29:0] core_io_ptw_pmp_4_addr; // @[RocketTile.scala 115:20]
  wire [31:0] core_io_ptw_pmp_4_mask; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_5_cfg_l; // @[RocketTile.scala 115:20]
  wire [1:0] core_io_ptw_pmp_5_cfg_a; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_5_cfg_x; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_5_cfg_w; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_5_cfg_r; // @[RocketTile.scala 115:20]
  wire [29:0] core_io_ptw_pmp_5_addr; // @[RocketTile.scala 115:20]
  wire [31:0] core_io_ptw_pmp_5_mask; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_6_cfg_l; // @[RocketTile.scala 115:20]
  wire [1:0] core_io_ptw_pmp_6_cfg_a; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_6_cfg_x; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_6_cfg_w; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_6_cfg_r; // @[RocketTile.scala 115:20]
  wire [29:0] core_io_ptw_pmp_6_addr; // @[RocketTile.scala 115:20]
  wire [31:0] core_io_ptw_pmp_6_mask; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_7_cfg_l; // @[RocketTile.scala 115:20]
  wire [1:0] core_io_ptw_pmp_7_cfg_a; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_7_cfg_x; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_7_cfg_w; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pmp_7_cfg_r; // @[RocketTile.scala 115:20]
  wire [29:0] core_io_ptw_pmp_7_addr; // @[RocketTile.scala 115:20]
  wire [31:0] core_io_ptw_pmp_7_mask; // @[RocketTile.scala 115:20]
  wire [63:0] core_io_ptw_customCSRs_csrs_0_value; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pcode_req_valid; // @[RocketTile.scala 115:20]
  wire [1:0] core_io_ptw_pcode_req_bits_id; // @[RocketTile.scala 115:20]
  wire [19:0] core_io_ptw_pcode_req_bits_value_base; // @[RocketTile.scala 115:20]
  wire [9:0] core_io_ptw_pcode_req_bits_value_mask; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pcode_req_bits_value_valid; // @[RocketTile.scala 115:20]
  wire  core_io_ptw_pcode_req_bits_value_locked; // @[RocketTile.scala 115:20]
  wire [26:0] core_io_ptw_vpoffset_req_bits_value; // @[RocketTile.scala 115:20]
  wire [31:0] core_io_fpu_inst; // @[RocketTile.scala 115:20]
  wire [63:0] core_io_fpu_fromint_data; // @[RocketTile.scala 115:20]
  wire [2:0] core_io_fpu_fcsr_rm; // @[RocketTile.scala 115:20]
  wire  core_io_fpu_fcsr_flags_valid; // @[RocketTile.scala 115:20]
  wire [4:0] core_io_fpu_fcsr_flags_bits; // @[RocketTile.scala 115:20]
  wire [63:0] core_io_fpu_store_data; // @[RocketTile.scala 115:20]
  wire [63:0] core_io_fpu_toint_data; // @[RocketTile.scala 115:20]
  wire  core_io_fpu_dmem_resp_val; // @[RocketTile.scala 115:20]
  wire [2:0] core_io_fpu_dmem_resp_type; // @[RocketTile.scala 115:20]
  wire [4:0] core_io_fpu_dmem_resp_tag; // @[RocketTile.scala 115:20]
  wire [63:0] core_io_fpu_dmem_resp_data; // @[RocketTile.scala 115:20]
  wire  core_io_fpu_valid; // @[RocketTile.scala 115:20]
  wire  core_io_fpu_fcsr_rdy; // @[RocketTile.scala 115:20]
  wire  core_io_fpu_nack_mem; // @[RocketTile.scala 115:20]
  wire  core_io_fpu_illegal_rm; // @[RocketTile.scala 115:20]
  wire  core_io_fpu_killx; // @[RocketTile.scala 115:20]
  wire  core_io_fpu_killm; // @[RocketTile.scala 115:20]
  wire  core_io_fpu_dec_wen; // @[RocketTile.scala 115:20]
  wire  core_io_fpu_dec_ren1; // @[RocketTile.scala 115:20]
  wire  core_io_fpu_dec_ren2; // @[RocketTile.scala 115:20]
  wire  core_io_fpu_dec_ren3; // @[RocketTile.scala 115:20]
  wire  core_io_fpu_sboard_set; // @[RocketTile.scala 115:20]
  wire  core_io_fpu_sboard_clr; // @[RocketTile.scala 115:20]
  wire [4:0] core_io_fpu_sboard_clra; // @[RocketTile.scala 115:20]
  wire [29:0] core_io_covSum; // @[RocketTile.scala 115:20]
  wire  core_metaAssert; // @[RocketTile.scala 115:20]
  wire  core_metaReset; // @[RocketTile.scala 115:20]
  wire  core_csr_halt; // @[RocketTile.scala 115:20]
  wire  core_div_halt; // @[RocketTile.scala 115:20]
  wire  core_ibuf_halt; // @[RocketTile.scala 115:20]
  wire [29:0] RocketTile_covSum;
  wire [29:0] intsink_1_sum;
  wire [29:0] intsink_sum;
  wire [29:0] dcache_sum;
  wire [29:0] dcacheArb_sum;
  wire [29:0] intsink_2_sum;
  wire [29:0] frontend_sum;
  wire [29:0] buffer_sum;
  wire [29:0] core_sum;
  wire [29:0] intsink_3_sum;
  wire [29:0] ptw_sum;
  wire [29:0] tlMasterXbar_sum;
  wire [29:0] fpuOpt_sum;
  wire [29:0] intXbar_sum;
  wire  ptw_metaAssert_wire;
  wire  intsink_2_metaAssert_wire;
  wire  intsink_metaAssert_wire;
  wire  fpuOpt_metaAssert_wire;
  wire  frontend_metaAssert_wire;
  wire  dcacheArb_metaAssert_wire;
  wire  buffer_metaAssert_wire;
  wire  intsink_1_metaAssert_wire;
  wire  intXbar_metaAssert_wire;
  wire  core_metaAssert_wire;
  wire  tlMasterXbar_metaAssert_wire;
  wire  intsink_3_metaAssert_wire;
  wire  dcache_metaAssert_wire;
  wire  RocketTile_or8;
  wire  RocketTile_or3;
  wire  RocketTile_or10;
  wire  RocketTile_or4;
  wire  RocketTile_or1;
  wire  RocketTile_or12;
  wire  RocketTile_or5;
  wire  RocketTile_or13;
  wire  RocketTile_or14;
  wire  RocketTile_or6;
  wire  RocketTile_or2;
  wire  RocketTile_or0;
  reg  RocketTile_metaAssert;
  reg [31:0] _RAND_0;
  TLXbar_8 tlMasterXbar ( // @[BaseTile.scala 142:42]
    .clock(tlMasterXbar_clock),
    .reset(tlMasterXbar_reset),
    .auto_in_1_a_ready(tlMasterXbar_auto_in_1_a_ready),
    .auto_in_1_a_valid(tlMasterXbar_auto_in_1_a_valid),
    .auto_in_1_a_bits_address(tlMasterXbar_auto_in_1_a_bits_address),
    .auto_in_1_d_valid(tlMasterXbar_auto_in_1_d_valid),
    .auto_in_1_d_bits_opcode(tlMasterXbar_auto_in_1_d_bits_opcode),
    .auto_in_1_d_bits_size(tlMasterXbar_auto_in_1_d_bits_size),
    .auto_in_1_d_bits_data(tlMasterXbar_auto_in_1_d_bits_data),
    .auto_in_1_d_bits_corrupt(tlMasterXbar_auto_in_1_d_bits_corrupt),
    .auto_in_0_a_ready(tlMasterXbar_auto_in_0_a_ready),
    .auto_in_0_a_valid(tlMasterXbar_auto_in_0_a_valid),
    .auto_in_0_a_bits_opcode(tlMasterXbar_auto_in_0_a_bits_opcode),
    .auto_in_0_a_bits_param(tlMasterXbar_auto_in_0_a_bits_param),
    .auto_in_0_a_bits_size(tlMasterXbar_auto_in_0_a_bits_size),
    .auto_in_0_a_bits_source(tlMasterXbar_auto_in_0_a_bits_source),
    .auto_in_0_a_bits_address(tlMasterXbar_auto_in_0_a_bits_address),
    .auto_in_0_a_bits_mask(tlMasterXbar_auto_in_0_a_bits_mask),
    .auto_in_0_a_bits_data(tlMasterXbar_auto_in_0_a_bits_data),
    .auto_in_0_b_ready(tlMasterXbar_auto_in_0_b_ready),
    .auto_in_0_b_valid(tlMasterXbar_auto_in_0_b_valid),
    .auto_in_0_b_bits_param(tlMasterXbar_auto_in_0_b_bits_param),
    .auto_in_0_b_bits_size(tlMasterXbar_auto_in_0_b_bits_size),
    .auto_in_0_b_bits_source(tlMasterXbar_auto_in_0_b_bits_source),
    .auto_in_0_b_bits_address(tlMasterXbar_auto_in_0_b_bits_address),
    .auto_in_0_c_ready(tlMasterXbar_auto_in_0_c_ready),
    .auto_in_0_c_valid(tlMasterXbar_auto_in_0_c_valid),
    .auto_in_0_c_bits_opcode(tlMasterXbar_auto_in_0_c_bits_opcode),
    .auto_in_0_c_bits_param(tlMasterXbar_auto_in_0_c_bits_param),
    .auto_in_0_c_bits_size(tlMasterXbar_auto_in_0_c_bits_size),
    .auto_in_0_c_bits_source(tlMasterXbar_auto_in_0_c_bits_source),
    .auto_in_0_c_bits_address(tlMasterXbar_auto_in_0_c_bits_address),
    .auto_in_0_c_bits_data(tlMasterXbar_auto_in_0_c_bits_data),
    .auto_in_0_d_ready(tlMasterXbar_auto_in_0_d_ready),
    .auto_in_0_d_valid(tlMasterXbar_auto_in_0_d_valid),
    .auto_in_0_d_bits_opcode(tlMasterXbar_auto_in_0_d_bits_opcode),
    .auto_in_0_d_bits_param(tlMasterXbar_auto_in_0_d_bits_param),
    .auto_in_0_d_bits_size(tlMasterXbar_auto_in_0_d_bits_size),
    .auto_in_0_d_bits_source(tlMasterXbar_auto_in_0_d_bits_source),
    .auto_in_0_d_bits_sink(tlMasterXbar_auto_in_0_d_bits_sink),
    .auto_in_0_d_bits_denied(tlMasterXbar_auto_in_0_d_bits_denied),
    .auto_in_0_d_bits_data(tlMasterXbar_auto_in_0_d_bits_data),
    .auto_in_0_e_ready(tlMasterXbar_auto_in_0_e_ready),
    .auto_in_0_e_valid(tlMasterXbar_auto_in_0_e_valid),
    .auto_in_0_e_bits_sink(tlMasterXbar_auto_in_0_e_bits_sink),
    .auto_out_a_ready(tlMasterXbar_auto_out_a_ready),
    .auto_out_a_valid(tlMasterXbar_auto_out_a_valid),
    .auto_out_a_bits_opcode(tlMasterXbar_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(tlMasterXbar_auto_out_a_bits_param),
    .auto_out_a_bits_size(tlMasterXbar_auto_out_a_bits_size),
    .auto_out_a_bits_source(tlMasterXbar_auto_out_a_bits_source),
    .auto_out_a_bits_address(tlMasterXbar_auto_out_a_bits_address),
    .auto_out_a_bits_mask(tlMasterXbar_auto_out_a_bits_mask),
    .auto_out_a_bits_data(tlMasterXbar_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(tlMasterXbar_auto_out_a_bits_corrupt),
    .auto_out_b_ready(tlMasterXbar_auto_out_b_ready),
    .auto_out_b_valid(tlMasterXbar_auto_out_b_valid),
    .auto_out_b_bits_opcode(tlMasterXbar_auto_out_b_bits_opcode),
    .auto_out_b_bits_param(tlMasterXbar_auto_out_b_bits_param),
    .auto_out_b_bits_size(tlMasterXbar_auto_out_b_bits_size),
    .auto_out_b_bits_source(tlMasterXbar_auto_out_b_bits_source),
    .auto_out_b_bits_address(tlMasterXbar_auto_out_b_bits_address),
    .auto_out_b_bits_mask(tlMasterXbar_auto_out_b_bits_mask),
    .auto_out_b_bits_corrupt(tlMasterXbar_auto_out_b_bits_corrupt),
    .auto_out_c_ready(tlMasterXbar_auto_out_c_ready),
    .auto_out_c_valid(tlMasterXbar_auto_out_c_valid),
    .auto_out_c_bits_opcode(tlMasterXbar_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(tlMasterXbar_auto_out_c_bits_param),
    .auto_out_c_bits_size(tlMasterXbar_auto_out_c_bits_size),
    .auto_out_c_bits_source(tlMasterXbar_auto_out_c_bits_source),
    .auto_out_c_bits_address(tlMasterXbar_auto_out_c_bits_address),
    .auto_out_c_bits_data(tlMasterXbar_auto_out_c_bits_data),
    .auto_out_d_ready(tlMasterXbar_auto_out_d_ready),
    .auto_out_d_valid(tlMasterXbar_auto_out_d_valid),
    .auto_out_d_bits_opcode(tlMasterXbar_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(tlMasterXbar_auto_out_d_bits_param),
    .auto_out_d_bits_size(tlMasterXbar_auto_out_d_bits_size),
    .auto_out_d_bits_source(tlMasterXbar_auto_out_d_bits_source),
    .auto_out_d_bits_sink(tlMasterXbar_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(tlMasterXbar_auto_out_d_bits_denied),
    .auto_out_d_bits_data(tlMasterXbar_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(tlMasterXbar_auto_out_d_bits_corrupt),
    .auto_out_e_ready(tlMasterXbar_auto_out_e_ready),
    .auto_out_e_valid(tlMasterXbar_auto_out_e_valid),
    .auto_out_e_bits_sink(tlMasterXbar_auto_out_e_bits_sink),
    .io_covSum(tlMasterXbar_io_covSum),
    .metaAssert(tlMasterXbar_metaAssert),
    .metaReset(tlMasterXbar_metaReset),
    .TLMonitor_halt(tlMasterXbar_TLMonitor_halt),
    .TLMonitor_1_halt(tlMasterXbar_TLMonitor_1_halt)
  );
  IntXbar_1 intXbar ( // @[BaseTile.scala 144:37]
    .auto_int_in_3_0(intXbar_auto_int_in_3_0),
    .auto_int_in_2_0(intXbar_auto_int_in_2_0),
    .auto_int_in_1_0(intXbar_auto_int_in_1_0),
    .auto_int_in_1_1(intXbar_auto_int_in_1_1),
    .auto_int_in_0_0(intXbar_auto_int_in_0_0),
    .auto_int_out_0(intXbar_auto_int_out_0),
    .auto_int_out_1(intXbar_auto_int_out_1),
    .auto_int_out_2(intXbar_auto_int_out_2),
    .auto_int_out_3(intXbar_auto_int_out_3),
    .auto_int_out_4(intXbar_auto_int_out_4),
    .io_covSum(intXbar_io_covSum),
    .metaAssert(intXbar_metaAssert)
  );
  DCache dcache ( // @[HellaCache.scala 215:43]
    .gated_clock(dcache_gated_clock),
    .reset(dcache_reset),
    .auto_out_a_ready(dcache_auto_out_a_ready),
    .auto_out_a_valid(dcache_auto_out_a_valid),
    .auto_out_a_bits_opcode(dcache_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(dcache_auto_out_a_bits_param),
    .auto_out_a_bits_size(dcache_auto_out_a_bits_size),
    .auto_out_a_bits_source(dcache_auto_out_a_bits_source),
    .auto_out_a_bits_address(dcache_auto_out_a_bits_address),
    .auto_out_a_bits_mask(dcache_auto_out_a_bits_mask),
    .auto_out_a_bits_data(dcache_auto_out_a_bits_data),
    .auto_out_b_ready(dcache_auto_out_b_ready),
    .auto_out_b_valid(dcache_auto_out_b_valid),
    .auto_out_b_bits_param(dcache_auto_out_b_bits_param),
    .auto_out_b_bits_size(dcache_auto_out_b_bits_size),
    .auto_out_b_bits_source(dcache_auto_out_b_bits_source),
    .auto_out_b_bits_address(dcache_auto_out_b_bits_address),
    .auto_out_c_ready(dcache_auto_out_c_ready),
    .auto_out_c_valid(dcache_auto_out_c_valid),
    .auto_out_c_bits_opcode(dcache_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(dcache_auto_out_c_bits_param),
    .auto_out_c_bits_size(dcache_auto_out_c_bits_size),
    .auto_out_c_bits_source(dcache_auto_out_c_bits_source),
    .auto_out_c_bits_address(dcache_auto_out_c_bits_address),
    .auto_out_c_bits_data(dcache_auto_out_c_bits_data),
    .auto_out_d_ready(dcache_auto_out_d_ready),
    .auto_out_d_valid(dcache_auto_out_d_valid),
    .auto_out_d_bits_opcode(dcache_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(dcache_auto_out_d_bits_param),
    .auto_out_d_bits_size(dcache_auto_out_d_bits_size),
    .auto_out_d_bits_source(dcache_auto_out_d_bits_source),
    .auto_out_d_bits_sink(dcache_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(dcache_auto_out_d_bits_denied),
    .auto_out_d_bits_data(dcache_auto_out_d_bits_data),
    .auto_out_e_ready(dcache_auto_out_e_ready),
    .auto_out_e_valid(dcache_auto_out_e_valid),
    .auto_out_e_bits_sink(dcache_auto_out_e_bits_sink),
    .io_cpu_req_ready(dcache_io_cpu_req_ready),
    .io_cpu_req_valid(dcache_io_cpu_req_valid),
    .io_cpu_req_bits_addr(dcache_io_cpu_req_bits_addr),
    .io_cpu_req_bits_tag(dcache_io_cpu_req_bits_tag),
    .io_cpu_req_bits_cmd(dcache_io_cpu_req_bits_cmd),
    .io_cpu_req_bits_typ(dcache_io_cpu_req_bits_typ),
    .io_cpu_req_bits_phys(dcache_io_cpu_req_bits_phys),
    .io_cpu_s1_kill(dcache_io_cpu_s1_kill),
    .io_cpu_s1_data_data(dcache_io_cpu_s1_data_data),
    .io_cpu_s2_nack(dcache_io_cpu_s2_nack),
    .io_cpu_resp_valid(dcache_io_cpu_resp_valid),
    .io_cpu_resp_bits_tag(dcache_io_cpu_resp_bits_tag),
    .io_cpu_resp_bits_typ(dcache_io_cpu_resp_bits_typ),
    .io_cpu_resp_bits_data(dcache_io_cpu_resp_bits_data),
    .io_cpu_resp_bits_replay(dcache_io_cpu_resp_bits_replay),
    .io_cpu_resp_bits_has_data(dcache_io_cpu_resp_bits_has_data),
    .io_cpu_resp_bits_data_word_bypass(dcache_io_cpu_resp_bits_data_word_bypass),
    .io_cpu_replay_next(dcache_io_cpu_replay_next),
    .io_cpu_s2_xcpt_ma_ld(dcache_io_cpu_s2_xcpt_ma_ld),
    .io_cpu_s2_xcpt_ma_st(dcache_io_cpu_s2_xcpt_ma_st),
    .io_cpu_s2_xcpt_pf_ld(dcache_io_cpu_s2_xcpt_pf_ld),
    .io_cpu_s2_xcpt_pf_st(dcache_io_cpu_s2_xcpt_pf_st),
    .io_cpu_s2_xcpt_ae_ld(dcache_io_cpu_s2_xcpt_ae_ld),
    .io_cpu_s2_xcpt_ae_st(dcache_io_cpu_s2_xcpt_ae_st),
    .io_cpu_ordered(dcache_io_cpu_ordered),
    .io_cpu_perf_grant(dcache_io_cpu_perf_grant),
    .io_cpu_keep_clock_enabled(dcache_io_cpu_keep_clock_enabled),
    .io_cpu_clock_enabled(dcache_io_cpu_clock_enabled),
    .io_ptw_req_ready(dcache_io_ptw_req_ready),
    .io_ptw_req_valid(dcache_io_ptw_req_valid),
    .io_ptw_req_bits_bits_addr(dcache_io_ptw_req_bits_bits_addr),
    .io_ptw_resp_valid(dcache_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae(dcache_io_ptw_resp_bits_ae),
    .io_ptw_resp_bits_pte_ppn(dcache_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d(dcache_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(dcache_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(dcache_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(dcache_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(dcache_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(dcache_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(dcache_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(dcache_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(dcache_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous(dcache_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(dcache_io_ptw_ptbr_mode),
    .io_ptw_status_dprv(dcache_io_ptw_status_dprv),
    .io_ptw_status_mxr(dcache_io_ptw_status_mxr),
    .io_ptw_status_sum(dcache_io_ptw_status_sum),
    .io_ptw_pmp_0_cfg_l(dcache_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a(dcache_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(dcache_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(dcache_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(dcache_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(dcache_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(dcache_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(dcache_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a(dcache_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(dcache_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(dcache_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(dcache_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(dcache_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(dcache_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(dcache_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a(dcache_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(dcache_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(dcache_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(dcache_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(dcache_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(dcache_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(dcache_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a(dcache_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(dcache_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(dcache_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(dcache_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(dcache_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(dcache_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(dcache_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a(dcache_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(dcache_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(dcache_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(dcache_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(dcache_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(dcache_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(dcache_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a(dcache_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(dcache_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(dcache_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(dcache_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(dcache_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(dcache_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(dcache_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a(dcache_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(dcache_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(dcache_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(dcache_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(dcache_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(dcache_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(dcache_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a(dcache_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(dcache_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(dcache_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(dcache_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(dcache_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(dcache_io_ptw_pmp_7_mask),
    .io_ptw_vpoffset_bits_value(dcache_io_ptw_vpoffset_bits_value),
    .io_covSum(dcache_io_covSum),
    .metaAssert(dcache_metaAssert),
    .metaReset(dcache_metaReset),
    .data_halt(dcache_data_halt),
    .tlb_halt(dcache_tlb_halt)
  );
  Frontend frontend ( // @[Frontend.scala 340:28]
    .gated_clock(frontend_gated_clock),
    .reset(frontend_reset),
    .auto_icache_master_out_a_ready(frontend_auto_icache_master_out_a_ready),
    .auto_icache_master_out_a_valid(frontend_auto_icache_master_out_a_valid),
    .auto_icache_master_out_a_bits_address(frontend_auto_icache_master_out_a_bits_address),
    .auto_icache_master_out_d_valid(frontend_auto_icache_master_out_d_valid),
    .auto_icache_master_out_d_bits_opcode(frontend_auto_icache_master_out_d_bits_opcode),
    .auto_icache_master_out_d_bits_size(frontend_auto_icache_master_out_d_bits_size),
    .auto_icache_master_out_d_bits_data(frontend_auto_icache_master_out_d_bits_data),
    .auto_icache_master_out_d_bits_corrupt(frontend_auto_icache_master_out_d_bits_corrupt),
    .io_reset_vector(frontend_io_reset_vector),
    .io_cpu_might_request(frontend_io_cpu_might_request),
    .io_cpu_req_valid(frontend_io_cpu_req_valid),
    .io_cpu_req_bits_pc(frontend_io_cpu_req_bits_pc),
    .io_cpu_req_bits_speculative(frontend_io_cpu_req_bits_speculative),
    .io_cpu_sfence_valid(frontend_io_cpu_sfence_valid),
    .io_cpu_sfence_bits_rs1(frontend_io_cpu_sfence_bits_rs1),
    .io_cpu_sfence_bits_rs2(frontend_io_cpu_sfence_bits_rs2),
    .io_cpu_sfence_bits_addr(frontend_io_cpu_sfence_bits_addr),
    .io_cpu_resp_ready(frontend_io_cpu_resp_ready),
    .io_cpu_resp_valid(frontend_io_cpu_resp_valid),
    .io_cpu_resp_bits_btb_taken(frontend_io_cpu_resp_bits_btb_taken),
    .io_cpu_resp_bits_btb_bridx(frontend_io_cpu_resp_bits_btb_bridx),
    .io_cpu_resp_bits_btb_entry(frontend_io_cpu_resp_bits_btb_entry),
    .io_cpu_resp_bits_btb_bht_history(frontend_io_cpu_resp_bits_btb_bht_history),
    .io_cpu_resp_bits_pc(frontend_io_cpu_resp_bits_pc),
    .io_cpu_resp_bits_data(frontend_io_cpu_resp_bits_data),
    .io_cpu_resp_bits_xcpt_pf_inst(frontend_io_cpu_resp_bits_xcpt_pf_inst),
    .io_cpu_resp_bits_xcpt_ae_inst(frontend_io_cpu_resp_bits_xcpt_ae_inst),
    .io_cpu_resp_bits_replay(frontend_io_cpu_resp_bits_replay),
    .io_cpu_btb_update_valid(frontend_io_cpu_btb_update_valid),
    .io_cpu_btb_update_bits_prediction_entry(frontend_io_cpu_btb_update_bits_prediction_entry),
    .io_cpu_btb_update_bits_pc(frontend_io_cpu_btb_update_bits_pc),
    .io_cpu_btb_update_bits_isValid(frontend_io_cpu_btb_update_bits_isValid),
    .io_cpu_btb_update_bits_br_pc(frontend_io_cpu_btb_update_bits_br_pc),
    .io_cpu_btb_update_bits_cfiType(frontend_io_cpu_btb_update_bits_cfiType),
    .io_cpu_bht_update_valid(frontend_io_cpu_bht_update_valid),
    .io_cpu_bht_update_bits_prediction_history(frontend_io_cpu_bht_update_bits_prediction_history),
    .io_cpu_bht_update_bits_pc(frontend_io_cpu_bht_update_bits_pc),
    .io_cpu_bht_update_bits_branch(frontend_io_cpu_bht_update_bits_branch),
    .io_cpu_bht_update_bits_taken(frontend_io_cpu_bht_update_bits_taken),
    .io_cpu_bht_update_bits_mispredict(frontend_io_cpu_bht_update_bits_mispredict),
    .io_cpu_flush_icache(frontend_io_cpu_flush_icache),
    .io_cpu_npc(frontend_io_cpu_npc),
    .io_ptw_req_ready(frontend_io_ptw_req_ready),
    .io_ptw_req_valid(frontend_io_ptw_req_valid),
    .io_ptw_req_bits_valid(frontend_io_ptw_req_bits_valid),
    .io_ptw_req_bits_bits_addr(frontend_io_ptw_req_bits_bits_addr),
    .io_ptw_resp_valid(frontend_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae(frontend_io_ptw_resp_bits_ae),
    .io_ptw_resp_bits_pte_ppn(frontend_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d(frontend_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(frontend_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(frontend_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(frontend_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(frontend_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(frontend_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(frontend_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(frontend_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(frontend_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous(frontend_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(frontend_io_ptw_ptbr_mode),
    .io_ptw_status_prv(frontend_io_ptw_status_prv),
    .io_ptw_pmp_0_cfg_l(frontend_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a(frontend_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(frontend_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(frontend_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(frontend_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(frontend_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(frontend_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(frontend_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a(frontend_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(frontend_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(frontend_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(frontend_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(frontend_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(frontend_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(frontend_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a(frontend_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(frontend_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(frontend_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(frontend_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(frontend_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(frontend_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(frontend_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a(frontend_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(frontend_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(frontend_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(frontend_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(frontend_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(frontend_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(frontend_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a(frontend_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(frontend_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(frontend_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(frontend_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(frontend_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(frontend_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(frontend_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a(frontend_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(frontend_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(frontend_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(frontend_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(frontend_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(frontend_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(frontend_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a(frontend_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(frontend_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(frontend_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(frontend_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(frontend_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(frontend_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(frontend_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a(frontend_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(frontend_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(frontend_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(frontend_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(frontend_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(frontend_io_ptw_pmp_7_mask),
    .io_ptw_vpoffset_bits_value(frontend_io_ptw_vpoffset_bits_value),
    .io_covSum(frontend_io_covSum),
    .metaAssert(frontend_metaAssert),
    .metaReset(frontend_metaReset),
    .icache_halt(frontend_icache_halt),
    .fq_halt(frontend_fq_halt),
    .tlb_halt(frontend_tlb_halt),
    .btb_halt(frontend_btb_halt)
  );
  TLBuffer_22 buffer ( // @[Buffer.scala 69:28]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_in_a_ready(buffer_auto_in_a_ready),
    .auto_in_a_valid(buffer_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(buffer_auto_in_a_bits_param),
    .auto_in_a_bits_size(buffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(buffer_auto_in_a_bits_source),
    .auto_in_a_bits_address(buffer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(buffer_auto_in_a_bits_corrupt),
    .auto_in_b_ready(buffer_auto_in_b_ready),
    .auto_in_b_valid(buffer_auto_in_b_valid),
    .auto_in_b_bits_opcode(buffer_auto_in_b_bits_opcode),
    .auto_in_b_bits_param(buffer_auto_in_b_bits_param),
    .auto_in_b_bits_size(buffer_auto_in_b_bits_size),
    .auto_in_b_bits_source(buffer_auto_in_b_bits_source),
    .auto_in_b_bits_address(buffer_auto_in_b_bits_address),
    .auto_in_b_bits_mask(buffer_auto_in_b_bits_mask),
    .auto_in_b_bits_corrupt(buffer_auto_in_b_bits_corrupt),
    .auto_in_c_ready(buffer_auto_in_c_ready),
    .auto_in_c_valid(buffer_auto_in_c_valid),
    .auto_in_c_bits_opcode(buffer_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(buffer_auto_in_c_bits_param),
    .auto_in_c_bits_size(buffer_auto_in_c_bits_size),
    .auto_in_c_bits_source(buffer_auto_in_c_bits_source),
    .auto_in_c_bits_address(buffer_auto_in_c_bits_address),
    .auto_in_c_bits_data(buffer_auto_in_c_bits_data),
    .auto_in_d_ready(buffer_auto_in_d_ready),
    .auto_in_d_valid(buffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(buffer_auto_in_d_bits_param),
    .auto_in_d_bits_size(buffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(buffer_auto_in_d_bits_source),
    .auto_in_d_bits_sink(buffer_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(buffer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
    .auto_in_e_ready(buffer_auto_in_e_ready),
    .auto_in_e_valid(buffer_auto_in_e_valid),
    .auto_in_e_bits_sink(buffer_auto_in_e_bits_sink),
    .auto_out_a_ready(buffer_auto_out_a_ready),
    .auto_out_a_valid(buffer_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(buffer_auto_out_a_bits_param),
    .auto_out_a_bits_size(buffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(buffer_auto_out_a_bits_corrupt),
    .auto_out_b_ready(buffer_auto_out_b_ready),
    .auto_out_b_valid(buffer_auto_out_b_valid),
    .auto_out_b_bits_opcode(buffer_auto_out_b_bits_opcode),
    .auto_out_b_bits_param(buffer_auto_out_b_bits_param),
    .auto_out_b_bits_size(buffer_auto_out_b_bits_size),
    .auto_out_b_bits_source(buffer_auto_out_b_bits_source),
    .auto_out_b_bits_address(buffer_auto_out_b_bits_address),
    .auto_out_b_bits_mask(buffer_auto_out_b_bits_mask),
    .auto_out_b_bits_corrupt(buffer_auto_out_b_bits_corrupt),
    .auto_out_c_ready(buffer_auto_out_c_ready),
    .auto_out_c_valid(buffer_auto_out_c_valid),
    .auto_out_c_bits_opcode(buffer_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(buffer_auto_out_c_bits_param),
    .auto_out_c_bits_size(buffer_auto_out_c_bits_size),
    .auto_out_c_bits_source(buffer_auto_out_c_bits_source),
    .auto_out_c_bits_address(buffer_auto_out_c_bits_address),
    .auto_out_c_bits_data(buffer_auto_out_c_bits_data),
    .auto_out_c_bits_corrupt(buffer_auto_out_c_bits_corrupt),
    .auto_out_d_ready(buffer_auto_out_d_ready),
    .auto_out_d_valid(buffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(buffer_auto_out_d_bits_param),
    .auto_out_d_bits_size(buffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_auto_out_d_bits_source),
    .auto_out_d_bits_sink(buffer_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(buffer_auto_out_d_bits_denied),
    .auto_out_d_bits_data(buffer_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(buffer_auto_out_d_bits_corrupt),
    .auto_out_e_ready(buffer_auto_out_e_ready),
    .auto_out_e_valid(buffer_auto_out_e_valid),
    .auto_out_e_bits_sink(buffer_auto_out_e_bits_sink),
    .io_covSum(buffer_io_covSum),
    .metaAssert(buffer_metaAssert),
    .metaReset(buffer_metaReset),
    .TLMonitor_halt(buffer_TLMonitor_halt),
    .Queue_4_halt(buffer_Queue_4_halt),
    .Queue_2_halt(buffer_Queue_2_halt),
    .Queue_1_halt(buffer_Queue_1_halt),
    .Queue_3_halt(buffer_Queue_3_halt),
    .Queue_halt(buffer_Queue_halt)
  );
  IntSyncCrossingSink intsink ( // @[Crossing.scala 63:29]
    .clock(intsink_clock),
    .auto_in_sync_0(intsink_auto_in_sync_0),
    .auto_out_0(intsink_auto_out_0),
    .io_covSum(intsink_io_covSum),
    .metaAssert(intsink_metaAssert),
    .metaReset(intsink_metaReset),
    .SynchronizerShiftReg_w1_d3_halt(intsink_SynchronizerShiftReg_w1_d3_halt)
  );
  IntSyncCrossingSink_1 intsink_1 ( // @[Crossing.scala 63:29]
    .auto_in_sync_0(intsink_1_auto_in_sync_0),
    .auto_in_sync_1(intsink_1_auto_in_sync_1),
    .auto_out_0(intsink_1_auto_out_0),
    .auto_out_1(intsink_1_auto_out_1),
    .io_covSum(intsink_1_io_covSum),
    .metaAssert(intsink_1_metaAssert)
  );
  IntSyncCrossingSink_2 intsink_2 ( // @[Crossing.scala 63:29]
    .auto_in_sync_0(intsink_2_auto_in_sync_0),
    .auto_out_0(intsink_2_auto_out_0),
    .io_covSum(intsink_2_io_covSum),
    .metaAssert(intsink_2_metaAssert)
  );
  IntSyncCrossingSink_2 intsink_3 ( // @[Crossing.scala 63:29]
    .auto_in_sync_0(intsink_3_auto_in_sync_0),
    .auto_out_0(intsink_3_auto_out_0),
    .io_covSum(intsink_3_io_covSum),
    .metaAssert(intsink_3_metaAssert)
  );
  FPU fpuOpt ( // @[RocketTile.scala 173:62]
    .clock(fpuOpt_clock),
    .reset(fpuOpt_reset),
    .io_inst(fpuOpt_io_inst),
    .io_fromint_data(fpuOpt_io_fromint_data),
    .io_fcsr_rm(fpuOpt_io_fcsr_rm),
    .io_fcsr_flags_valid(fpuOpt_io_fcsr_flags_valid),
    .io_fcsr_flags_bits(fpuOpt_io_fcsr_flags_bits),
    .io_store_data(fpuOpt_io_store_data),
    .io_toint_data(fpuOpt_io_toint_data),
    .io_dmem_resp_val(fpuOpt_io_dmem_resp_val),
    .io_dmem_resp_type(fpuOpt_io_dmem_resp_type),
    .io_dmem_resp_tag(fpuOpt_io_dmem_resp_tag),
    .io_dmem_resp_data(fpuOpt_io_dmem_resp_data),
    .io_valid(fpuOpt_io_valid),
    .io_fcsr_rdy(fpuOpt_io_fcsr_rdy),
    .io_nack_mem(fpuOpt_io_nack_mem),
    .io_illegal_rm(fpuOpt_io_illegal_rm),
    .io_killx(fpuOpt_io_killx),
    .io_killm(fpuOpt_io_killm),
    .io_dec_wen(fpuOpt_io_dec_wen),
    .io_dec_ren1(fpuOpt_io_dec_ren1),
    .io_dec_ren2(fpuOpt_io_dec_ren2),
    .io_dec_ren3(fpuOpt_io_dec_ren3),
    .io_sboard_set(fpuOpt_io_sboard_set),
    .io_sboard_clr(fpuOpt_io_sboard_clr),
    .io_sboard_clra(fpuOpt_io_sboard_clra),
    .io_covSum(fpuOpt_io_covSum),
    .metaAssert(fpuOpt_metaAssert),
    .metaReset(fpuOpt_metaReset),
    .dfma_halt(fpuOpt_dfma_halt),
    .fpmu_halt(fpuOpt_fpmu_halt),
    .divSqrt_1_halt(fpuOpt_divSqrt_1_halt),
    .ifpu_halt(fpuOpt_ifpu_halt),
    .divSqrt_halt(fpuOpt_divSqrt_halt),
    .fpiu_halt(fpuOpt_fpiu_halt),
    .sfma_halt(fpuOpt_sfma_halt)
  );
  HellaCacheArbiter dcacheArb ( // @[HellaCache.scala 227:25]
    .clock(dcacheArb_clock),
    .io_requestor_0_req_ready(dcacheArb_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(dcacheArb_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_addr(dcacheArb_io_requestor_0_req_bits_addr),
    .io_requestor_0_s1_kill(dcacheArb_io_requestor_0_s1_kill),
    .io_requestor_0_s2_nack(dcacheArb_io_requestor_0_s2_nack),
    .io_requestor_0_resp_valid(dcacheArb_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_data_word_bypass(dcacheArb_io_requestor_0_resp_bits_data_word_bypass),
    .io_requestor_0_s2_xcpt_ae_ld(dcacheArb_io_requestor_0_s2_xcpt_ae_ld),
    .io_requestor_1_req_ready(dcacheArb_io_requestor_1_req_ready),
    .io_requestor_1_req_valid(dcacheArb_io_requestor_1_req_valid),
    .io_requestor_1_req_bits_addr(dcacheArb_io_requestor_1_req_bits_addr),
    .io_requestor_1_req_bits_tag(dcacheArb_io_requestor_1_req_bits_tag),
    .io_requestor_1_req_bits_cmd(dcacheArb_io_requestor_1_req_bits_cmd),
    .io_requestor_1_req_bits_typ(dcacheArb_io_requestor_1_req_bits_typ),
    .io_requestor_1_s1_kill(dcacheArb_io_requestor_1_s1_kill),
    .io_requestor_1_s1_data_data(dcacheArb_io_requestor_1_s1_data_data),
    .io_requestor_1_s2_nack(dcacheArb_io_requestor_1_s2_nack),
    .io_requestor_1_resp_valid(dcacheArb_io_requestor_1_resp_valid),
    .io_requestor_1_resp_bits_tag(dcacheArb_io_requestor_1_resp_bits_tag),
    .io_requestor_1_resp_bits_typ(dcacheArb_io_requestor_1_resp_bits_typ),
    .io_requestor_1_resp_bits_data(dcacheArb_io_requestor_1_resp_bits_data),
    .io_requestor_1_resp_bits_replay(dcacheArb_io_requestor_1_resp_bits_replay),
    .io_requestor_1_resp_bits_has_data(dcacheArb_io_requestor_1_resp_bits_has_data),
    .io_requestor_1_resp_bits_data_word_bypass(dcacheArb_io_requestor_1_resp_bits_data_word_bypass),
    .io_requestor_1_replay_next(dcacheArb_io_requestor_1_replay_next),
    .io_requestor_1_s2_xcpt_ma_ld(dcacheArb_io_requestor_1_s2_xcpt_ma_ld),
    .io_requestor_1_s2_xcpt_ma_st(dcacheArb_io_requestor_1_s2_xcpt_ma_st),
    .io_requestor_1_s2_xcpt_pf_ld(dcacheArb_io_requestor_1_s2_xcpt_pf_ld),
    .io_requestor_1_s2_xcpt_pf_st(dcacheArb_io_requestor_1_s2_xcpt_pf_st),
    .io_requestor_1_s2_xcpt_ae_ld(dcacheArb_io_requestor_1_s2_xcpt_ae_ld),
    .io_requestor_1_s2_xcpt_ae_st(dcacheArb_io_requestor_1_s2_xcpt_ae_st),
    .io_requestor_1_ordered(dcacheArb_io_requestor_1_ordered),
    .io_requestor_1_perf_grant(dcacheArb_io_requestor_1_perf_grant),
    .io_requestor_1_keep_clock_enabled(dcacheArb_io_requestor_1_keep_clock_enabled),
    .io_requestor_1_clock_enabled(dcacheArb_io_requestor_1_clock_enabled),
    .io_mem_req_ready(dcacheArb_io_mem_req_ready),
    .io_mem_req_valid(dcacheArb_io_mem_req_valid),
    .io_mem_req_bits_addr(dcacheArb_io_mem_req_bits_addr),
    .io_mem_req_bits_tag(dcacheArb_io_mem_req_bits_tag),
    .io_mem_req_bits_cmd(dcacheArb_io_mem_req_bits_cmd),
    .io_mem_req_bits_typ(dcacheArb_io_mem_req_bits_typ),
    .io_mem_req_bits_phys(dcacheArb_io_mem_req_bits_phys),
    .io_mem_s1_kill(dcacheArb_io_mem_s1_kill),
    .io_mem_s1_data_data(dcacheArb_io_mem_s1_data_data),
    .io_mem_s2_nack(dcacheArb_io_mem_s2_nack),
    .io_mem_resp_valid(dcacheArb_io_mem_resp_valid),
    .io_mem_resp_bits_tag(dcacheArb_io_mem_resp_bits_tag),
    .io_mem_resp_bits_typ(dcacheArb_io_mem_resp_bits_typ),
    .io_mem_resp_bits_data(dcacheArb_io_mem_resp_bits_data),
    .io_mem_resp_bits_replay(dcacheArb_io_mem_resp_bits_replay),
    .io_mem_resp_bits_has_data(dcacheArb_io_mem_resp_bits_has_data),
    .io_mem_resp_bits_data_word_bypass(dcacheArb_io_mem_resp_bits_data_word_bypass),
    .io_mem_replay_next(dcacheArb_io_mem_replay_next),
    .io_mem_s2_xcpt_ma_ld(dcacheArb_io_mem_s2_xcpt_ma_ld),
    .io_mem_s2_xcpt_ma_st(dcacheArb_io_mem_s2_xcpt_ma_st),
    .io_mem_s2_xcpt_pf_ld(dcacheArb_io_mem_s2_xcpt_pf_ld),
    .io_mem_s2_xcpt_pf_st(dcacheArb_io_mem_s2_xcpt_pf_st),
    .io_mem_s2_xcpt_ae_ld(dcacheArb_io_mem_s2_xcpt_ae_ld),
    .io_mem_s2_xcpt_ae_st(dcacheArb_io_mem_s2_xcpt_ae_st),
    .io_mem_ordered(dcacheArb_io_mem_ordered),
    .io_mem_perf_grant(dcacheArb_io_mem_perf_grant),
    .io_mem_keep_clock_enabled(dcacheArb_io_mem_keep_clock_enabled),
    .io_mem_clock_enabled(dcacheArb_io_mem_clock_enabled),
    .io_covSum(dcacheArb_io_covSum),
    .metaAssert(dcacheArb_metaAssert),
    .metaReset(dcacheArb_metaReset)
  );
  PTW ptw ( // @[PTW.scala 531:19]
    .clock(ptw_clock),
    .reset(ptw_reset),
    .io_requestor_0_req_ready(ptw_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(ptw_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_bits_addr(ptw_io_requestor_0_req_bits_bits_addr),
    .io_requestor_0_resp_valid(ptw_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_ae(ptw_io_requestor_0_resp_bits_ae),
    .io_requestor_0_resp_bits_pte_ppn(ptw_io_requestor_0_resp_bits_pte_ppn),
    .io_requestor_0_resp_bits_pte_d(ptw_io_requestor_0_resp_bits_pte_d),
    .io_requestor_0_resp_bits_pte_a(ptw_io_requestor_0_resp_bits_pte_a),
    .io_requestor_0_resp_bits_pte_g(ptw_io_requestor_0_resp_bits_pte_g),
    .io_requestor_0_resp_bits_pte_u(ptw_io_requestor_0_resp_bits_pte_u),
    .io_requestor_0_resp_bits_pte_x(ptw_io_requestor_0_resp_bits_pte_x),
    .io_requestor_0_resp_bits_pte_w(ptw_io_requestor_0_resp_bits_pte_w),
    .io_requestor_0_resp_bits_pte_r(ptw_io_requestor_0_resp_bits_pte_r),
    .io_requestor_0_resp_bits_pte_v(ptw_io_requestor_0_resp_bits_pte_v),
    .io_requestor_0_resp_bits_level(ptw_io_requestor_0_resp_bits_level),
    .io_requestor_0_resp_bits_homogeneous(ptw_io_requestor_0_resp_bits_homogeneous),
    .io_requestor_0_ptbr_mode(ptw_io_requestor_0_ptbr_mode),
    .io_requestor_0_status_dprv(ptw_io_requestor_0_status_dprv),
    .io_requestor_0_status_mxr(ptw_io_requestor_0_status_mxr),
    .io_requestor_0_status_sum(ptw_io_requestor_0_status_sum),
    .io_requestor_0_pmp_0_cfg_l(ptw_io_requestor_0_pmp_0_cfg_l),
    .io_requestor_0_pmp_0_cfg_a(ptw_io_requestor_0_pmp_0_cfg_a),
    .io_requestor_0_pmp_0_cfg_x(ptw_io_requestor_0_pmp_0_cfg_x),
    .io_requestor_0_pmp_0_cfg_w(ptw_io_requestor_0_pmp_0_cfg_w),
    .io_requestor_0_pmp_0_cfg_r(ptw_io_requestor_0_pmp_0_cfg_r),
    .io_requestor_0_pmp_0_addr(ptw_io_requestor_0_pmp_0_addr),
    .io_requestor_0_pmp_0_mask(ptw_io_requestor_0_pmp_0_mask),
    .io_requestor_0_pmp_1_cfg_l(ptw_io_requestor_0_pmp_1_cfg_l),
    .io_requestor_0_pmp_1_cfg_a(ptw_io_requestor_0_pmp_1_cfg_a),
    .io_requestor_0_pmp_1_cfg_x(ptw_io_requestor_0_pmp_1_cfg_x),
    .io_requestor_0_pmp_1_cfg_w(ptw_io_requestor_0_pmp_1_cfg_w),
    .io_requestor_0_pmp_1_cfg_r(ptw_io_requestor_0_pmp_1_cfg_r),
    .io_requestor_0_pmp_1_addr(ptw_io_requestor_0_pmp_1_addr),
    .io_requestor_0_pmp_1_mask(ptw_io_requestor_0_pmp_1_mask),
    .io_requestor_0_pmp_2_cfg_l(ptw_io_requestor_0_pmp_2_cfg_l),
    .io_requestor_0_pmp_2_cfg_a(ptw_io_requestor_0_pmp_2_cfg_a),
    .io_requestor_0_pmp_2_cfg_x(ptw_io_requestor_0_pmp_2_cfg_x),
    .io_requestor_0_pmp_2_cfg_w(ptw_io_requestor_0_pmp_2_cfg_w),
    .io_requestor_0_pmp_2_cfg_r(ptw_io_requestor_0_pmp_2_cfg_r),
    .io_requestor_0_pmp_2_addr(ptw_io_requestor_0_pmp_2_addr),
    .io_requestor_0_pmp_2_mask(ptw_io_requestor_0_pmp_2_mask),
    .io_requestor_0_pmp_3_cfg_l(ptw_io_requestor_0_pmp_3_cfg_l),
    .io_requestor_0_pmp_3_cfg_a(ptw_io_requestor_0_pmp_3_cfg_a),
    .io_requestor_0_pmp_3_cfg_x(ptw_io_requestor_0_pmp_3_cfg_x),
    .io_requestor_0_pmp_3_cfg_w(ptw_io_requestor_0_pmp_3_cfg_w),
    .io_requestor_0_pmp_3_cfg_r(ptw_io_requestor_0_pmp_3_cfg_r),
    .io_requestor_0_pmp_3_addr(ptw_io_requestor_0_pmp_3_addr),
    .io_requestor_0_pmp_3_mask(ptw_io_requestor_0_pmp_3_mask),
    .io_requestor_0_pmp_4_cfg_l(ptw_io_requestor_0_pmp_4_cfg_l),
    .io_requestor_0_pmp_4_cfg_a(ptw_io_requestor_0_pmp_4_cfg_a),
    .io_requestor_0_pmp_4_cfg_x(ptw_io_requestor_0_pmp_4_cfg_x),
    .io_requestor_0_pmp_4_cfg_w(ptw_io_requestor_0_pmp_4_cfg_w),
    .io_requestor_0_pmp_4_cfg_r(ptw_io_requestor_0_pmp_4_cfg_r),
    .io_requestor_0_pmp_4_addr(ptw_io_requestor_0_pmp_4_addr),
    .io_requestor_0_pmp_4_mask(ptw_io_requestor_0_pmp_4_mask),
    .io_requestor_0_pmp_5_cfg_l(ptw_io_requestor_0_pmp_5_cfg_l),
    .io_requestor_0_pmp_5_cfg_a(ptw_io_requestor_0_pmp_5_cfg_a),
    .io_requestor_0_pmp_5_cfg_x(ptw_io_requestor_0_pmp_5_cfg_x),
    .io_requestor_0_pmp_5_cfg_w(ptw_io_requestor_0_pmp_5_cfg_w),
    .io_requestor_0_pmp_5_cfg_r(ptw_io_requestor_0_pmp_5_cfg_r),
    .io_requestor_0_pmp_5_addr(ptw_io_requestor_0_pmp_5_addr),
    .io_requestor_0_pmp_5_mask(ptw_io_requestor_0_pmp_5_mask),
    .io_requestor_0_pmp_6_cfg_l(ptw_io_requestor_0_pmp_6_cfg_l),
    .io_requestor_0_pmp_6_cfg_a(ptw_io_requestor_0_pmp_6_cfg_a),
    .io_requestor_0_pmp_6_cfg_x(ptw_io_requestor_0_pmp_6_cfg_x),
    .io_requestor_0_pmp_6_cfg_w(ptw_io_requestor_0_pmp_6_cfg_w),
    .io_requestor_0_pmp_6_cfg_r(ptw_io_requestor_0_pmp_6_cfg_r),
    .io_requestor_0_pmp_6_addr(ptw_io_requestor_0_pmp_6_addr),
    .io_requestor_0_pmp_6_mask(ptw_io_requestor_0_pmp_6_mask),
    .io_requestor_0_pmp_7_cfg_l(ptw_io_requestor_0_pmp_7_cfg_l),
    .io_requestor_0_pmp_7_cfg_a(ptw_io_requestor_0_pmp_7_cfg_a),
    .io_requestor_0_pmp_7_cfg_x(ptw_io_requestor_0_pmp_7_cfg_x),
    .io_requestor_0_pmp_7_cfg_w(ptw_io_requestor_0_pmp_7_cfg_w),
    .io_requestor_0_pmp_7_cfg_r(ptw_io_requestor_0_pmp_7_cfg_r),
    .io_requestor_0_pmp_7_addr(ptw_io_requestor_0_pmp_7_addr),
    .io_requestor_0_pmp_7_mask(ptw_io_requestor_0_pmp_7_mask),
    .io_requestor_0_vpoffset_bits_value(ptw_io_requestor_0_vpoffset_bits_value),
    .io_requestor_1_req_ready(ptw_io_requestor_1_req_ready),
    .io_requestor_1_req_valid(ptw_io_requestor_1_req_valid),
    .io_requestor_1_req_bits_valid(ptw_io_requestor_1_req_bits_valid),
    .io_requestor_1_req_bits_bits_addr(ptw_io_requestor_1_req_bits_bits_addr),
    .io_requestor_1_resp_valid(ptw_io_requestor_1_resp_valid),
    .io_requestor_1_resp_bits_ae(ptw_io_requestor_1_resp_bits_ae),
    .io_requestor_1_resp_bits_pte_ppn(ptw_io_requestor_1_resp_bits_pte_ppn),
    .io_requestor_1_resp_bits_pte_d(ptw_io_requestor_1_resp_bits_pte_d),
    .io_requestor_1_resp_bits_pte_a(ptw_io_requestor_1_resp_bits_pte_a),
    .io_requestor_1_resp_bits_pte_g(ptw_io_requestor_1_resp_bits_pte_g),
    .io_requestor_1_resp_bits_pte_u(ptw_io_requestor_1_resp_bits_pte_u),
    .io_requestor_1_resp_bits_pte_x(ptw_io_requestor_1_resp_bits_pte_x),
    .io_requestor_1_resp_bits_pte_w(ptw_io_requestor_1_resp_bits_pte_w),
    .io_requestor_1_resp_bits_pte_r(ptw_io_requestor_1_resp_bits_pte_r),
    .io_requestor_1_resp_bits_pte_v(ptw_io_requestor_1_resp_bits_pte_v),
    .io_requestor_1_resp_bits_level(ptw_io_requestor_1_resp_bits_level),
    .io_requestor_1_resp_bits_homogeneous(ptw_io_requestor_1_resp_bits_homogeneous),
    .io_requestor_1_ptbr_mode(ptw_io_requestor_1_ptbr_mode),
    .io_requestor_1_status_prv(ptw_io_requestor_1_status_prv),
    .io_requestor_1_pmp_0_cfg_l(ptw_io_requestor_1_pmp_0_cfg_l),
    .io_requestor_1_pmp_0_cfg_a(ptw_io_requestor_1_pmp_0_cfg_a),
    .io_requestor_1_pmp_0_cfg_x(ptw_io_requestor_1_pmp_0_cfg_x),
    .io_requestor_1_pmp_0_cfg_w(ptw_io_requestor_1_pmp_0_cfg_w),
    .io_requestor_1_pmp_0_cfg_r(ptw_io_requestor_1_pmp_0_cfg_r),
    .io_requestor_1_pmp_0_addr(ptw_io_requestor_1_pmp_0_addr),
    .io_requestor_1_pmp_0_mask(ptw_io_requestor_1_pmp_0_mask),
    .io_requestor_1_pmp_1_cfg_l(ptw_io_requestor_1_pmp_1_cfg_l),
    .io_requestor_1_pmp_1_cfg_a(ptw_io_requestor_1_pmp_1_cfg_a),
    .io_requestor_1_pmp_1_cfg_x(ptw_io_requestor_1_pmp_1_cfg_x),
    .io_requestor_1_pmp_1_cfg_w(ptw_io_requestor_1_pmp_1_cfg_w),
    .io_requestor_1_pmp_1_cfg_r(ptw_io_requestor_1_pmp_1_cfg_r),
    .io_requestor_1_pmp_1_addr(ptw_io_requestor_1_pmp_1_addr),
    .io_requestor_1_pmp_1_mask(ptw_io_requestor_1_pmp_1_mask),
    .io_requestor_1_pmp_2_cfg_l(ptw_io_requestor_1_pmp_2_cfg_l),
    .io_requestor_1_pmp_2_cfg_a(ptw_io_requestor_1_pmp_2_cfg_a),
    .io_requestor_1_pmp_2_cfg_x(ptw_io_requestor_1_pmp_2_cfg_x),
    .io_requestor_1_pmp_2_cfg_w(ptw_io_requestor_1_pmp_2_cfg_w),
    .io_requestor_1_pmp_2_cfg_r(ptw_io_requestor_1_pmp_2_cfg_r),
    .io_requestor_1_pmp_2_addr(ptw_io_requestor_1_pmp_2_addr),
    .io_requestor_1_pmp_2_mask(ptw_io_requestor_1_pmp_2_mask),
    .io_requestor_1_pmp_3_cfg_l(ptw_io_requestor_1_pmp_3_cfg_l),
    .io_requestor_1_pmp_3_cfg_a(ptw_io_requestor_1_pmp_3_cfg_a),
    .io_requestor_1_pmp_3_cfg_x(ptw_io_requestor_1_pmp_3_cfg_x),
    .io_requestor_1_pmp_3_cfg_w(ptw_io_requestor_1_pmp_3_cfg_w),
    .io_requestor_1_pmp_3_cfg_r(ptw_io_requestor_1_pmp_3_cfg_r),
    .io_requestor_1_pmp_3_addr(ptw_io_requestor_1_pmp_3_addr),
    .io_requestor_1_pmp_3_mask(ptw_io_requestor_1_pmp_3_mask),
    .io_requestor_1_pmp_4_cfg_l(ptw_io_requestor_1_pmp_4_cfg_l),
    .io_requestor_1_pmp_4_cfg_a(ptw_io_requestor_1_pmp_4_cfg_a),
    .io_requestor_1_pmp_4_cfg_x(ptw_io_requestor_1_pmp_4_cfg_x),
    .io_requestor_1_pmp_4_cfg_w(ptw_io_requestor_1_pmp_4_cfg_w),
    .io_requestor_1_pmp_4_cfg_r(ptw_io_requestor_1_pmp_4_cfg_r),
    .io_requestor_1_pmp_4_addr(ptw_io_requestor_1_pmp_4_addr),
    .io_requestor_1_pmp_4_mask(ptw_io_requestor_1_pmp_4_mask),
    .io_requestor_1_pmp_5_cfg_l(ptw_io_requestor_1_pmp_5_cfg_l),
    .io_requestor_1_pmp_5_cfg_a(ptw_io_requestor_1_pmp_5_cfg_a),
    .io_requestor_1_pmp_5_cfg_x(ptw_io_requestor_1_pmp_5_cfg_x),
    .io_requestor_1_pmp_5_cfg_w(ptw_io_requestor_1_pmp_5_cfg_w),
    .io_requestor_1_pmp_5_cfg_r(ptw_io_requestor_1_pmp_5_cfg_r),
    .io_requestor_1_pmp_5_addr(ptw_io_requestor_1_pmp_5_addr),
    .io_requestor_1_pmp_5_mask(ptw_io_requestor_1_pmp_5_mask),
    .io_requestor_1_pmp_6_cfg_l(ptw_io_requestor_1_pmp_6_cfg_l),
    .io_requestor_1_pmp_6_cfg_a(ptw_io_requestor_1_pmp_6_cfg_a),
    .io_requestor_1_pmp_6_cfg_x(ptw_io_requestor_1_pmp_6_cfg_x),
    .io_requestor_1_pmp_6_cfg_w(ptw_io_requestor_1_pmp_6_cfg_w),
    .io_requestor_1_pmp_6_cfg_r(ptw_io_requestor_1_pmp_6_cfg_r),
    .io_requestor_1_pmp_6_addr(ptw_io_requestor_1_pmp_6_addr),
    .io_requestor_1_pmp_6_mask(ptw_io_requestor_1_pmp_6_mask),
    .io_requestor_1_pmp_7_cfg_l(ptw_io_requestor_1_pmp_7_cfg_l),
    .io_requestor_1_pmp_7_cfg_a(ptw_io_requestor_1_pmp_7_cfg_a),
    .io_requestor_1_pmp_7_cfg_x(ptw_io_requestor_1_pmp_7_cfg_x),
    .io_requestor_1_pmp_7_cfg_w(ptw_io_requestor_1_pmp_7_cfg_w),
    .io_requestor_1_pmp_7_cfg_r(ptw_io_requestor_1_pmp_7_cfg_r),
    .io_requestor_1_pmp_7_addr(ptw_io_requestor_1_pmp_7_addr),
    .io_requestor_1_pmp_7_mask(ptw_io_requestor_1_pmp_7_mask),
    .io_requestor_1_vpoffset_bits_value(ptw_io_requestor_1_vpoffset_bits_value),
    .io_mem_req_ready(ptw_io_mem_req_ready),
    .io_mem_req_valid(ptw_io_mem_req_valid),
    .io_mem_req_bits_addr(ptw_io_mem_req_bits_addr),
    .io_mem_s1_kill(ptw_io_mem_s1_kill),
    .io_mem_s2_nack(ptw_io_mem_s2_nack),
    .io_mem_resp_valid(ptw_io_mem_resp_valid),
    .io_mem_resp_bits_data_word_bypass(ptw_io_mem_resp_bits_data_word_bypass),
    .io_mem_s2_xcpt_ae_ld(ptw_io_mem_s2_xcpt_ae_ld),
    .io_dpath_ptbr_mode(ptw_io_dpath_ptbr_mode),
    .io_dpath_ptbr_ppn(ptw_io_dpath_ptbr_ppn),
    .io_dpath_sfence_valid(ptw_io_dpath_sfence_valid),
    .io_dpath_sfence_bits_rs1(ptw_io_dpath_sfence_bits_rs1),
    .io_dpath_status_dprv(ptw_io_dpath_status_dprv),
    .io_dpath_status_prv(ptw_io_dpath_status_prv),
    .io_dpath_status_mxr(ptw_io_dpath_status_mxr),
    .io_dpath_status_sum(ptw_io_dpath_status_sum),
    .io_dpath_pmp_0_cfg_l(ptw_io_dpath_pmp_0_cfg_l),
    .io_dpath_pmp_0_cfg_a(ptw_io_dpath_pmp_0_cfg_a),
    .io_dpath_pmp_0_cfg_x(ptw_io_dpath_pmp_0_cfg_x),
    .io_dpath_pmp_0_cfg_w(ptw_io_dpath_pmp_0_cfg_w),
    .io_dpath_pmp_0_cfg_r(ptw_io_dpath_pmp_0_cfg_r),
    .io_dpath_pmp_0_addr(ptw_io_dpath_pmp_0_addr),
    .io_dpath_pmp_0_mask(ptw_io_dpath_pmp_0_mask),
    .io_dpath_pmp_1_cfg_l(ptw_io_dpath_pmp_1_cfg_l),
    .io_dpath_pmp_1_cfg_a(ptw_io_dpath_pmp_1_cfg_a),
    .io_dpath_pmp_1_cfg_x(ptw_io_dpath_pmp_1_cfg_x),
    .io_dpath_pmp_1_cfg_w(ptw_io_dpath_pmp_1_cfg_w),
    .io_dpath_pmp_1_cfg_r(ptw_io_dpath_pmp_1_cfg_r),
    .io_dpath_pmp_1_addr(ptw_io_dpath_pmp_1_addr),
    .io_dpath_pmp_1_mask(ptw_io_dpath_pmp_1_mask),
    .io_dpath_pmp_2_cfg_l(ptw_io_dpath_pmp_2_cfg_l),
    .io_dpath_pmp_2_cfg_a(ptw_io_dpath_pmp_2_cfg_a),
    .io_dpath_pmp_2_cfg_x(ptw_io_dpath_pmp_2_cfg_x),
    .io_dpath_pmp_2_cfg_w(ptw_io_dpath_pmp_2_cfg_w),
    .io_dpath_pmp_2_cfg_r(ptw_io_dpath_pmp_2_cfg_r),
    .io_dpath_pmp_2_addr(ptw_io_dpath_pmp_2_addr),
    .io_dpath_pmp_2_mask(ptw_io_dpath_pmp_2_mask),
    .io_dpath_pmp_3_cfg_l(ptw_io_dpath_pmp_3_cfg_l),
    .io_dpath_pmp_3_cfg_a(ptw_io_dpath_pmp_3_cfg_a),
    .io_dpath_pmp_3_cfg_x(ptw_io_dpath_pmp_3_cfg_x),
    .io_dpath_pmp_3_cfg_w(ptw_io_dpath_pmp_3_cfg_w),
    .io_dpath_pmp_3_cfg_r(ptw_io_dpath_pmp_3_cfg_r),
    .io_dpath_pmp_3_addr(ptw_io_dpath_pmp_3_addr),
    .io_dpath_pmp_3_mask(ptw_io_dpath_pmp_3_mask),
    .io_dpath_pmp_4_cfg_l(ptw_io_dpath_pmp_4_cfg_l),
    .io_dpath_pmp_4_cfg_a(ptw_io_dpath_pmp_4_cfg_a),
    .io_dpath_pmp_4_cfg_x(ptw_io_dpath_pmp_4_cfg_x),
    .io_dpath_pmp_4_cfg_w(ptw_io_dpath_pmp_4_cfg_w),
    .io_dpath_pmp_4_cfg_r(ptw_io_dpath_pmp_4_cfg_r),
    .io_dpath_pmp_4_addr(ptw_io_dpath_pmp_4_addr),
    .io_dpath_pmp_4_mask(ptw_io_dpath_pmp_4_mask),
    .io_dpath_pmp_5_cfg_l(ptw_io_dpath_pmp_5_cfg_l),
    .io_dpath_pmp_5_cfg_a(ptw_io_dpath_pmp_5_cfg_a),
    .io_dpath_pmp_5_cfg_x(ptw_io_dpath_pmp_5_cfg_x),
    .io_dpath_pmp_5_cfg_w(ptw_io_dpath_pmp_5_cfg_w),
    .io_dpath_pmp_5_cfg_r(ptw_io_dpath_pmp_5_cfg_r),
    .io_dpath_pmp_5_addr(ptw_io_dpath_pmp_5_addr),
    .io_dpath_pmp_5_mask(ptw_io_dpath_pmp_5_mask),
    .io_dpath_pmp_6_cfg_l(ptw_io_dpath_pmp_6_cfg_l),
    .io_dpath_pmp_6_cfg_a(ptw_io_dpath_pmp_6_cfg_a),
    .io_dpath_pmp_6_cfg_x(ptw_io_dpath_pmp_6_cfg_x),
    .io_dpath_pmp_6_cfg_w(ptw_io_dpath_pmp_6_cfg_w),
    .io_dpath_pmp_6_cfg_r(ptw_io_dpath_pmp_6_cfg_r),
    .io_dpath_pmp_6_addr(ptw_io_dpath_pmp_6_addr),
    .io_dpath_pmp_6_mask(ptw_io_dpath_pmp_6_mask),
    .io_dpath_pmp_7_cfg_l(ptw_io_dpath_pmp_7_cfg_l),
    .io_dpath_pmp_7_cfg_a(ptw_io_dpath_pmp_7_cfg_a),
    .io_dpath_pmp_7_cfg_x(ptw_io_dpath_pmp_7_cfg_x),
    .io_dpath_pmp_7_cfg_w(ptw_io_dpath_pmp_7_cfg_w),
    .io_dpath_pmp_7_cfg_r(ptw_io_dpath_pmp_7_cfg_r),
    .io_dpath_pmp_7_addr(ptw_io_dpath_pmp_7_addr),
    .io_dpath_pmp_7_mask(ptw_io_dpath_pmp_7_mask),
    .io_dpath_pcode_req_valid(ptw_io_dpath_pcode_req_valid),
    .io_dpath_pcode_req_bits_id(ptw_io_dpath_pcode_req_bits_id),
    .io_dpath_pcode_req_bits_value_base(ptw_io_dpath_pcode_req_bits_value_base),
    .io_dpath_pcode_req_bits_value_mask(ptw_io_dpath_pcode_req_bits_value_mask),
    .io_dpath_pcode_req_bits_value_valid(ptw_io_dpath_pcode_req_bits_value_valid),
    .io_dpath_pcode_req_bits_value_locked(ptw_io_dpath_pcode_req_bits_value_locked),
    .io_dpath_vpoffset_req_bits_value(ptw_io_dpath_vpoffset_req_bits_value),
    .io_covSum(ptw_io_covSum),
    .metaAssert(ptw_metaAssert),
    .metaReset(ptw_metaReset),
    .arb_halt(ptw_arb_halt)
  );
  Rocket core ( // @[RocketTile.scala 115:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_hartid(core_io_hartid),
    .io_interrupts_debug(core_io_interrupts_debug),
    .io_interrupts_mtip(core_io_interrupts_mtip),
    .io_interrupts_msip(core_io_interrupts_msip),
    .io_interrupts_meip(core_io_interrupts_meip),
    .io_interrupts_seip(core_io_interrupts_seip),
    .io_imem_might_request(core_io_imem_might_request),
    .io_imem_req_valid(core_io_imem_req_valid),
    .io_imem_req_bits_pc(core_io_imem_req_bits_pc),
    .io_imem_req_bits_speculative(core_io_imem_req_bits_speculative),
    .io_imem_sfence_valid(core_io_imem_sfence_valid),
    .io_imem_sfence_bits_rs1(core_io_imem_sfence_bits_rs1),
    .io_imem_sfence_bits_rs2(core_io_imem_sfence_bits_rs2),
    .io_imem_sfence_bits_addr(core_io_imem_sfence_bits_addr),
    .io_imem_resp_ready(core_io_imem_resp_ready),
    .io_imem_resp_valid(core_io_imem_resp_valid),
    .io_imem_resp_bits_btb_taken(core_io_imem_resp_bits_btb_taken),
    .io_imem_resp_bits_btb_bridx(core_io_imem_resp_bits_btb_bridx),
    .io_imem_resp_bits_btb_entry(core_io_imem_resp_bits_btb_entry),
    .io_imem_resp_bits_btb_bht_history(core_io_imem_resp_bits_btb_bht_history),
    .io_imem_resp_bits_pc(core_io_imem_resp_bits_pc),
    .io_imem_resp_bits_data(core_io_imem_resp_bits_data),
    .io_imem_resp_bits_xcpt_pf_inst(core_io_imem_resp_bits_xcpt_pf_inst),
    .io_imem_resp_bits_xcpt_ae_inst(core_io_imem_resp_bits_xcpt_ae_inst),
    .io_imem_resp_bits_replay(core_io_imem_resp_bits_replay),
    .io_imem_btb_update_valid(core_io_imem_btb_update_valid),
    .io_imem_btb_update_bits_prediction_entry(core_io_imem_btb_update_bits_prediction_entry),
    .io_imem_btb_update_bits_pc(core_io_imem_btb_update_bits_pc),
    .io_imem_btb_update_bits_isValid(core_io_imem_btb_update_bits_isValid),
    .io_imem_btb_update_bits_br_pc(core_io_imem_btb_update_bits_br_pc),
    .io_imem_btb_update_bits_cfiType(core_io_imem_btb_update_bits_cfiType),
    .io_imem_bht_update_valid(core_io_imem_bht_update_valid),
    .io_imem_bht_update_bits_prediction_history(core_io_imem_bht_update_bits_prediction_history),
    .io_imem_bht_update_bits_pc(core_io_imem_bht_update_bits_pc),
    .io_imem_bht_update_bits_branch(core_io_imem_bht_update_bits_branch),
    .io_imem_bht_update_bits_taken(core_io_imem_bht_update_bits_taken),
    .io_imem_bht_update_bits_mispredict(core_io_imem_bht_update_bits_mispredict),
    .io_imem_flush_icache(core_io_imem_flush_icache),
    .io_dmem_req_ready(core_io_dmem_req_ready),
    .io_dmem_req_valid(core_io_dmem_req_valid),
    .io_dmem_req_bits_addr(core_io_dmem_req_bits_addr),
    .io_dmem_req_bits_tag(core_io_dmem_req_bits_tag),
    .io_dmem_req_bits_cmd(core_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_typ(core_io_dmem_req_bits_typ),
    .io_dmem_s1_kill(core_io_dmem_s1_kill),
    .io_dmem_s1_data_data(core_io_dmem_s1_data_data),
    .io_dmem_s2_nack(core_io_dmem_s2_nack),
    .io_dmem_resp_valid(core_io_dmem_resp_valid),
    .io_dmem_resp_bits_tag(core_io_dmem_resp_bits_tag),
    .io_dmem_resp_bits_typ(core_io_dmem_resp_bits_typ),
    .io_dmem_resp_bits_data(core_io_dmem_resp_bits_data),
    .io_dmem_resp_bits_replay(core_io_dmem_resp_bits_replay),
    .io_dmem_resp_bits_has_data(core_io_dmem_resp_bits_has_data),
    .io_dmem_resp_bits_data_word_bypass(core_io_dmem_resp_bits_data_word_bypass),
    .io_dmem_replay_next(core_io_dmem_replay_next),
    .io_dmem_s2_xcpt_ma_ld(core_io_dmem_s2_xcpt_ma_ld),
    .io_dmem_s2_xcpt_ma_st(core_io_dmem_s2_xcpt_ma_st),
    .io_dmem_s2_xcpt_pf_ld(core_io_dmem_s2_xcpt_pf_ld),
    .io_dmem_s2_xcpt_pf_st(core_io_dmem_s2_xcpt_pf_st),
    .io_dmem_s2_xcpt_ae_ld(core_io_dmem_s2_xcpt_ae_ld),
    .io_dmem_s2_xcpt_ae_st(core_io_dmem_s2_xcpt_ae_st),
    .io_dmem_ordered(core_io_dmem_ordered),
    .io_dmem_perf_grant(core_io_dmem_perf_grant),
    .io_dmem_keep_clock_enabled(core_io_dmem_keep_clock_enabled),
    .io_dmem_clock_enabled(core_io_dmem_clock_enabled),
    .io_ptw_ptbr_mode(core_io_ptw_ptbr_mode),
    .io_ptw_ptbr_ppn(core_io_ptw_ptbr_ppn),
    .io_ptw_sfence_valid(core_io_ptw_sfence_valid),
    .io_ptw_sfence_bits_rs1(core_io_ptw_sfence_bits_rs1),
    .io_ptw_status_dprv(core_io_ptw_status_dprv),
    .io_ptw_status_prv(core_io_ptw_status_prv),
    .io_ptw_status_mxr(core_io_ptw_status_mxr),
    .io_ptw_status_sum(core_io_ptw_status_sum),
    .io_ptw_pmp_0_cfg_l(core_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a(core_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(core_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(core_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(core_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(core_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(core_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(core_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a(core_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(core_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(core_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(core_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(core_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(core_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(core_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a(core_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(core_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(core_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(core_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(core_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(core_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(core_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a(core_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(core_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(core_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(core_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(core_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(core_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(core_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a(core_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(core_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(core_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(core_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(core_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(core_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(core_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a(core_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(core_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(core_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(core_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(core_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(core_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(core_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a(core_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(core_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(core_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(core_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(core_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(core_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(core_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a(core_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(core_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(core_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(core_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(core_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(core_io_ptw_pmp_7_mask),
    .io_ptw_customCSRs_csrs_0_value(core_io_ptw_customCSRs_csrs_0_value),
    .io_ptw_pcode_req_valid(core_io_ptw_pcode_req_valid),
    .io_ptw_pcode_req_bits_id(core_io_ptw_pcode_req_bits_id),
    .io_ptw_pcode_req_bits_value_base(core_io_ptw_pcode_req_bits_value_base),
    .io_ptw_pcode_req_bits_value_mask(core_io_ptw_pcode_req_bits_value_mask),
    .io_ptw_pcode_req_bits_value_valid(core_io_ptw_pcode_req_bits_value_valid),
    .io_ptw_pcode_req_bits_value_locked(core_io_ptw_pcode_req_bits_value_locked),
    .io_ptw_vpoffset_req_bits_value(core_io_ptw_vpoffset_req_bits_value),
    .io_fpu_inst(core_io_fpu_inst),
    .io_fpu_fromint_data(core_io_fpu_fromint_data),
    .io_fpu_fcsr_rm(core_io_fpu_fcsr_rm),
    .io_fpu_fcsr_flags_valid(core_io_fpu_fcsr_flags_valid),
    .io_fpu_fcsr_flags_bits(core_io_fpu_fcsr_flags_bits),
    .io_fpu_store_data(core_io_fpu_store_data),
    .io_fpu_toint_data(core_io_fpu_toint_data),
    .io_fpu_dmem_resp_val(core_io_fpu_dmem_resp_val),
    .io_fpu_dmem_resp_type(core_io_fpu_dmem_resp_type),
    .io_fpu_dmem_resp_tag(core_io_fpu_dmem_resp_tag),
    .io_fpu_dmem_resp_data(core_io_fpu_dmem_resp_data),
    .io_fpu_valid(core_io_fpu_valid),
    .io_fpu_fcsr_rdy(core_io_fpu_fcsr_rdy),
    .io_fpu_nack_mem(core_io_fpu_nack_mem),
    .io_fpu_illegal_rm(core_io_fpu_illegal_rm),
    .io_fpu_killx(core_io_fpu_killx),
    .io_fpu_killm(core_io_fpu_killm),
    .io_fpu_dec_wen(core_io_fpu_dec_wen),
    .io_fpu_dec_ren1(core_io_fpu_dec_ren1),
    .io_fpu_dec_ren2(core_io_fpu_dec_ren2),
    .io_fpu_dec_ren3(core_io_fpu_dec_ren3),
    .io_fpu_sboard_set(core_io_fpu_sboard_set),
    .io_fpu_sboard_clr(core_io_fpu_sboard_clr),
    .io_fpu_sboard_clra(core_io_fpu_sboard_clra),
    .io_covSum(core_io_covSum),
    .metaAssert(core_metaAssert),
    .metaReset(core_metaReset),
    .csr_halt(core_csr_halt),
    .div_halt(core_div_halt),
    .ibuf_halt(core_ibuf_halt)
  );
  assign auto_tl_master_xing_out_a_valid = buffer_auto_out_a_valid; // @[LazyModule.scala 173:49]
  assign auto_tl_master_xing_out_a_bits_opcode = buffer_auto_out_a_bits_opcode; // @[LazyModule.scala 173:49]
  assign auto_tl_master_xing_out_a_bits_param = buffer_auto_out_a_bits_param; // @[LazyModule.scala 173:49]
  assign auto_tl_master_xing_out_a_bits_size = buffer_auto_out_a_bits_size; // @[LazyModule.scala 173:49]
  assign auto_tl_master_xing_out_a_bits_source = buffer_auto_out_a_bits_source; // @[LazyModule.scala 173:49]
  assign auto_tl_master_xing_out_a_bits_address = buffer_auto_out_a_bits_address; // @[LazyModule.scala 173:49]
  assign auto_tl_master_xing_out_a_bits_mask = buffer_auto_out_a_bits_mask; // @[LazyModule.scala 173:49]
  assign auto_tl_master_xing_out_a_bits_data = buffer_auto_out_a_bits_data; // @[LazyModule.scala 173:49]
  assign auto_tl_master_xing_out_a_bits_corrupt = buffer_auto_out_a_bits_corrupt; // @[LazyModule.scala 173:49]
  assign auto_tl_master_xing_out_b_ready = buffer_auto_out_b_ready; // @[LazyModule.scala 173:49]
  assign auto_tl_master_xing_out_c_valid = buffer_auto_out_c_valid; // @[LazyModule.scala 173:49]
  assign auto_tl_master_xing_out_c_bits_opcode = buffer_auto_out_c_bits_opcode; // @[LazyModule.scala 173:49]
  assign auto_tl_master_xing_out_c_bits_param = buffer_auto_out_c_bits_param; // @[LazyModule.scala 173:49]
  assign auto_tl_master_xing_out_c_bits_size = buffer_auto_out_c_bits_size; // @[LazyModule.scala 173:49]
  assign auto_tl_master_xing_out_c_bits_source = buffer_auto_out_c_bits_source; // @[LazyModule.scala 173:49]
  assign auto_tl_master_xing_out_c_bits_address = buffer_auto_out_c_bits_address; // @[LazyModule.scala 173:49]
  assign auto_tl_master_xing_out_c_bits_data = buffer_auto_out_c_bits_data; // @[LazyModule.scala 173:49]
  assign auto_tl_master_xing_out_c_bits_corrupt = buffer_auto_out_c_bits_corrupt; // @[LazyModule.scala 173:49]
  assign auto_tl_master_xing_out_d_ready = buffer_auto_out_d_ready; // @[LazyModule.scala 173:49]
  assign auto_tl_master_xing_out_e_valid = buffer_auto_out_e_valid; // @[LazyModule.scala 173:49]
  assign auto_tl_master_xing_out_e_bits_sink = buffer_auto_out_e_bits_sink; // @[LazyModule.scala 173:49]
  assign tlMasterXbar_clock = clock;
  assign tlMasterXbar_reset = reset;
  assign tlMasterXbar_auto_in_1_a_valid = frontend_auto_icache_master_out_a_valid; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_in_1_a_bits_address = frontend_auto_icache_master_out_a_bits_address; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_in_0_a_valid = dcache_auto_out_a_valid; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_in_0_a_bits_opcode = dcache_auto_out_a_bits_opcode; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_in_0_a_bits_param = dcache_auto_out_a_bits_param; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_in_0_a_bits_size = dcache_auto_out_a_bits_size; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_in_0_a_bits_source = dcache_auto_out_a_bits_source; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_in_0_a_bits_address = dcache_auto_out_a_bits_address; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_in_0_a_bits_mask = dcache_auto_out_a_bits_mask; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_in_0_a_bits_data = dcache_auto_out_a_bits_data; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_in_0_b_ready = dcache_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_in_0_c_valid = dcache_auto_out_c_valid; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_in_0_c_bits_opcode = dcache_auto_out_c_bits_opcode; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_in_0_c_bits_param = dcache_auto_out_c_bits_param; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_in_0_c_bits_size = dcache_auto_out_c_bits_size; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_in_0_c_bits_source = dcache_auto_out_c_bits_source; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_in_0_c_bits_address = dcache_auto_out_c_bits_address; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_in_0_c_bits_data = dcache_auto_out_c_bits_data; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_in_0_d_ready = dcache_auto_out_d_ready; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_in_0_e_valid = dcache_auto_out_e_valid; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_in_0_e_bits_sink = dcache_auto_out_e_bits_sink; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_out_a_ready = buffer_auto_in_a_ready; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_out_b_valid = buffer_auto_in_b_valid; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_out_b_bits_opcode = buffer_auto_in_b_bits_opcode; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_out_b_bits_param = buffer_auto_in_b_bits_param; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_out_b_bits_size = buffer_auto_in_b_bits_size; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_out_b_bits_source = buffer_auto_in_b_bits_source; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_out_b_bits_address = buffer_auto_in_b_bits_address; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_out_b_bits_mask = buffer_auto_in_b_bits_mask; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_out_b_bits_corrupt = buffer_auto_in_b_bits_corrupt; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_out_c_ready = buffer_auto_in_c_ready; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_out_d_valid = buffer_auto_in_d_valid; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_out_d_bits_opcode = buffer_auto_in_d_bits_opcode; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_out_d_bits_param = buffer_auto_in_d_bits_param; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_out_d_bits_size = buffer_auto_in_d_bits_size; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_out_d_bits_source = buffer_auto_in_d_bits_source; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_out_d_bits_sink = buffer_auto_in_d_bits_sink; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_out_d_bits_denied = buffer_auto_in_d_bits_denied; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_out_d_bits_data = buffer_auto_in_d_bits_data; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_out_d_bits_corrupt = buffer_auto_in_d_bits_corrupt; // @[LazyModule.scala 167:31]
  assign tlMasterXbar_auto_out_e_ready = buffer_auto_in_e_ready; // @[LazyModule.scala 167:31]
  assign intXbar_auto_int_in_3_0 = intsink_3_auto_out_0; // @[LazyModule.scala 167:57]
  assign intXbar_auto_int_in_2_0 = intsink_2_auto_out_0; // @[LazyModule.scala 167:57]
  assign intXbar_auto_int_in_1_0 = intsink_1_auto_out_0; // @[LazyModule.scala 167:57]
  assign intXbar_auto_int_in_1_1 = intsink_1_auto_out_1; // @[LazyModule.scala 167:57]
  assign intXbar_auto_int_in_0_0 = intsink_auto_out_0; // @[LazyModule.scala 167:57]
  assign dcache_gated_clock = clock;
  assign dcache_reset = reset;
  assign dcache_auto_out_a_ready = tlMasterXbar_auto_in_0_a_ready; // @[LazyModule.scala 167:31]
  assign dcache_auto_out_b_valid = tlMasterXbar_auto_in_0_b_valid; // @[LazyModule.scala 167:31]
  assign dcache_auto_out_b_bits_param = tlMasterXbar_auto_in_0_b_bits_param; // @[LazyModule.scala 167:31]
  assign dcache_auto_out_b_bits_size = tlMasterXbar_auto_in_0_b_bits_size; // @[LazyModule.scala 167:31]
  assign dcache_auto_out_b_bits_source = tlMasterXbar_auto_in_0_b_bits_source; // @[LazyModule.scala 167:31]
  assign dcache_auto_out_b_bits_address = tlMasterXbar_auto_in_0_b_bits_address; // @[LazyModule.scala 167:31]
  assign dcache_auto_out_c_ready = tlMasterXbar_auto_in_0_c_ready; // @[LazyModule.scala 167:31]
  assign dcache_auto_out_d_valid = tlMasterXbar_auto_in_0_d_valid; // @[LazyModule.scala 167:31]
  assign dcache_auto_out_d_bits_opcode = tlMasterXbar_auto_in_0_d_bits_opcode; // @[LazyModule.scala 167:31]
  assign dcache_auto_out_d_bits_param = tlMasterXbar_auto_in_0_d_bits_param; // @[LazyModule.scala 167:31]
  assign dcache_auto_out_d_bits_size = tlMasterXbar_auto_in_0_d_bits_size; // @[LazyModule.scala 167:31]
  assign dcache_auto_out_d_bits_source = tlMasterXbar_auto_in_0_d_bits_source; // @[LazyModule.scala 167:31]
  assign dcache_auto_out_d_bits_sink = tlMasterXbar_auto_in_0_d_bits_sink; // @[LazyModule.scala 167:31]
  assign dcache_auto_out_d_bits_denied = tlMasterXbar_auto_in_0_d_bits_denied; // @[LazyModule.scala 167:31]
  assign dcache_auto_out_d_bits_data = tlMasterXbar_auto_in_0_d_bits_data; // @[LazyModule.scala 167:31]
  assign dcache_auto_out_e_ready = tlMasterXbar_auto_in_0_e_ready; // @[LazyModule.scala 167:31]
  assign dcache_io_cpu_req_valid = dcacheArb_io_mem_req_valid; // @[HellaCache.scala 228:30]
  assign dcache_io_cpu_req_bits_addr = dcacheArb_io_mem_req_bits_addr; // @[HellaCache.scala 228:30]
  assign dcache_io_cpu_req_bits_tag = dcacheArb_io_mem_req_bits_tag; // @[HellaCache.scala 228:30]
  assign dcache_io_cpu_req_bits_cmd = dcacheArb_io_mem_req_bits_cmd; // @[HellaCache.scala 228:30]
  assign dcache_io_cpu_req_bits_typ = dcacheArb_io_mem_req_bits_typ; // @[HellaCache.scala 228:30]
  assign dcache_io_cpu_req_bits_phys = dcacheArb_io_mem_req_bits_phys; // @[HellaCache.scala 228:30]
  assign dcache_io_cpu_s1_kill = dcacheArb_io_mem_s1_kill; // @[HellaCache.scala 228:30]
  assign dcache_io_cpu_s1_data_data = dcacheArb_io_mem_s1_data_data; // @[HellaCache.scala 228:30]
  assign dcache_io_cpu_keep_clock_enabled = dcacheArb_io_mem_keep_clock_enabled; // @[HellaCache.scala 228:30]
  assign dcache_io_ptw_req_ready = ptw_io_requestor_0_req_ready; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_resp_valid = ptw_io_requestor_0_resp_valid; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_resp_bits_ae = ptw_io_requestor_0_resp_bits_ae; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_resp_bits_pte_ppn = ptw_io_requestor_0_resp_bits_pte_ppn; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_resp_bits_pte_d = ptw_io_requestor_0_resp_bits_pte_d; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_resp_bits_pte_a = ptw_io_requestor_0_resp_bits_pte_a; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_resp_bits_pte_g = ptw_io_requestor_0_resp_bits_pte_g; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_resp_bits_pte_u = ptw_io_requestor_0_resp_bits_pte_u; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_resp_bits_pte_x = ptw_io_requestor_0_resp_bits_pte_x; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_resp_bits_pte_w = ptw_io_requestor_0_resp_bits_pte_w; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_resp_bits_pte_r = ptw_io_requestor_0_resp_bits_pte_r; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_resp_bits_pte_v = ptw_io_requestor_0_resp_bits_pte_v; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_resp_bits_level = ptw_io_requestor_0_resp_bits_level; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_resp_bits_homogeneous = ptw_io_requestor_0_resp_bits_homogeneous; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_ptbr_mode = ptw_io_requestor_0_ptbr_mode; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_status_dprv = ptw_io_requestor_0_status_dprv; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_status_mxr = ptw_io_requestor_0_status_mxr; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_status_sum = ptw_io_requestor_0_status_sum; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_0_cfg_l = ptw_io_requestor_0_pmp_0_cfg_l; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_0_cfg_a = ptw_io_requestor_0_pmp_0_cfg_a; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_0_cfg_x = ptw_io_requestor_0_pmp_0_cfg_x; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_0_cfg_w = ptw_io_requestor_0_pmp_0_cfg_w; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_0_cfg_r = ptw_io_requestor_0_pmp_0_cfg_r; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_0_addr = ptw_io_requestor_0_pmp_0_addr; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_0_mask = ptw_io_requestor_0_pmp_0_mask; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_1_cfg_l = ptw_io_requestor_0_pmp_1_cfg_l; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_1_cfg_a = ptw_io_requestor_0_pmp_1_cfg_a; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_1_cfg_x = ptw_io_requestor_0_pmp_1_cfg_x; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_1_cfg_w = ptw_io_requestor_0_pmp_1_cfg_w; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_1_cfg_r = ptw_io_requestor_0_pmp_1_cfg_r; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_1_addr = ptw_io_requestor_0_pmp_1_addr; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_1_mask = ptw_io_requestor_0_pmp_1_mask; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_2_cfg_l = ptw_io_requestor_0_pmp_2_cfg_l; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_2_cfg_a = ptw_io_requestor_0_pmp_2_cfg_a; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_2_cfg_x = ptw_io_requestor_0_pmp_2_cfg_x; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_2_cfg_w = ptw_io_requestor_0_pmp_2_cfg_w; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_2_cfg_r = ptw_io_requestor_0_pmp_2_cfg_r; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_2_addr = ptw_io_requestor_0_pmp_2_addr; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_2_mask = ptw_io_requestor_0_pmp_2_mask; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_3_cfg_l = ptw_io_requestor_0_pmp_3_cfg_l; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_3_cfg_a = ptw_io_requestor_0_pmp_3_cfg_a; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_3_cfg_x = ptw_io_requestor_0_pmp_3_cfg_x; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_3_cfg_w = ptw_io_requestor_0_pmp_3_cfg_w; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_3_cfg_r = ptw_io_requestor_0_pmp_3_cfg_r; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_3_addr = ptw_io_requestor_0_pmp_3_addr; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_3_mask = ptw_io_requestor_0_pmp_3_mask; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_4_cfg_l = ptw_io_requestor_0_pmp_4_cfg_l; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_4_cfg_a = ptw_io_requestor_0_pmp_4_cfg_a; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_4_cfg_x = ptw_io_requestor_0_pmp_4_cfg_x; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_4_cfg_w = ptw_io_requestor_0_pmp_4_cfg_w; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_4_cfg_r = ptw_io_requestor_0_pmp_4_cfg_r; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_4_addr = ptw_io_requestor_0_pmp_4_addr; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_4_mask = ptw_io_requestor_0_pmp_4_mask; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_5_cfg_l = ptw_io_requestor_0_pmp_5_cfg_l; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_5_cfg_a = ptw_io_requestor_0_pmp_5_cfg_a; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_5_cfg_x = ptw_io_requestor_0_pmp_5_cfg_x; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_5_cfg_w = ptw_io_requestor_0_pmp_5_cfg_w; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_5_cfg_r = ptw_io_requestor_0_pmp_5_cfg_r; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_5_addr = ptw_io_requestor_0_pmp_5_addr; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_5_mask = ptw_io_requestor_0_pmp_5_mask; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_6_cfg_l = ptw_io_requestor_0_pmp_6_cfg_l; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_6_cfg_a = ptw_io_requestor_0_pmp_6_cfg_a; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_6_cfg_x = ptw_io_requestor_0_pmp_6_cfg_x; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_6_cfg_w = ptw_io_requestor_0_pmp_6_cfg_w; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_6_cfg_r = ptw_io_requestor_0_pmp_6_cfg_r; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_6_addr = ptw_io_requestor_0_pmp_6_addr; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_6_mask = ptw_io_requestor_0_pmp_6_mask; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_7_cfg_l = ptw_io_requestor_0_pmp_7_cfg_l; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_7_cfg_a = ptw_io_requestor_0_pmp_7_cfg_a; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_7_cfg_x = ptw_io_requestor_0_pmp_7_cfg_x; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_7_cfg_w = ptw_io_requestor_0_pmp_7_cfg_w; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_7_cfg_r = ptw_io_requestor_0_pmp_7_cfg_r; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_7_addr = ptw_io_requestor_0_pmp_7_addr; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_pmp_7_mask = ptw_io_requestor_0_pmp_7_mask; // @[RocketTile.scala 169:20]
  assign dcache_io_ptw_vpoffset_bits_value = ptw_io_requestor_0_vpoffset_bits_value; // @[RocketTile.scala 169:20]
  assign frontend_gated_clock = clock;
  assign frontend_reset = reset;
  assign frontend_auto_icache_master_out_a_ready = tlMasterXbar_auto_in_1_a_ready; // @[LazyModule.scala 167:31]
  assign frontend_auto_icache_master_out_d_valid = tlMasterXbar_auto_in_1_d_valid; // @[LazyModule.scala 167:31]
  assign frontend_auto_icache_master_out_d_bits_opcode = tlMasterXbar_auto_in_1_d_bits_opcode; // @[LazyModule.scala 167:31]
  assign frontend_auto_icache_master_out_d_bits_size = tlMasterXbar_auto_in_1_d_bits_size; // @[LazyModule.scala 167:31]
  assign frontend_auto_icache_master_out_d_bits_data = tlMasterXbar_auto_in_1_d_bits_data; // @[LazyModule.scala 167:31]
  assign frontend_auto_icache_master_out_d_bits_corrupt = tlMasterXbar_auto_in_1_d_bits_corrupt; // @[LazyModule.scala 167:31]
  assign frontend_io_reset_vector = constants_reset_vector; // @[RocketTile.scala 131:41]
  assign frontend_io_cpu_might_request = core_io_imem_might_request; // @[RocketTile.scala 130:32]
  assign frontend_io_cpu_req_valid = core_io_imem_req_valid; // @[RocketTile.scala 130:32]
  assign frontend_io_cpu_req_bits_pc = core_io_imem_req_bits_pc; // @[RocketTile.scala 130:32]
  assign frontend_io_cpu_req_bits_speculative = core_io_imem_req_bits_speculative; // @[RocketTile.scala 130:32]
  assign frontend_io_cpu_sfence_valid = core_io_imem_sfence_valid; // @[RocketTile.scala 130:32]
  assign frontend_io_cpu_sfence_bits_rs1 = core_io_imem_sfence_bits_rs1; // @[RocketTile.scala 130:32]
  assign frontend_io_cpu_sfence_bits_rs2 = core_io_imem_sfence_bits_rs2; // @[RocketTile.scala 130:32]
  assign frontend_io_cpu_sfence_bits_addr = core_io_imem_sfence_bits_addr; // @[RocketTile.scala 130:32]
  assign frontend_io_cpu_resp_ready = core_io_imem_resp_ready; // @[RocketTile.scala 130:32]
  assign frontend_io_cpu_btb_update_valid = core_io_imem_btb_update_valid; // @[RocketTile.scala 130:32]
  assign frontend_io_cpu_btb_update_bits_prediction_entry = core_io_imem_btb_update_bits_prediction_entry; // @[RocketTile.scala 130:32]
  assign frontend_io_cpu_btb_update_bits_pc = core_io_imem_btb_update_bits_pc; // @[RocketTile.scala 130:32]
  assign frontend_io_cpu_btb_update_bits_isValid = core_io_imem_btb_update_bits_isValid; // @[RocketTile.scala 130:32]
  assign frontend_io_cpu_btb_update_bits_br_pc = core_io_imem_btb_update_bits_br_pc; // @[RocketTile.scala 130:32]
  assign frontend_io_cpu_btb_update_bits_cfiType = core_io_imem_btb_update_bits_cfiType; // @[RocketTile.scala 130:32]
  assign frontend_io_cpu_bht_update_valid = core_io_imem_bht_update_valid; // @[RocketTile.scala 130:32]
  assign frontend_io_cpu_bht_update_bits_prediction_history = core_io_imem_bht_update_bits_prediction_history; // @[RocketTile.scala 130:32]
  assign frontend_io_cpu_bht_update_bits_pc = core_io_imem_bht_update_bits_pc; // @[RocketTile.scala 130:32]
  assign frontend_io_cpu_bht_update_bits_branch = core_io_imem_bht_update_bits_branch; // @[RocketTile.scala 130:32]
  assign frontend_io_cpu_bht_update_bits_taken = core_io_imem_bht_update_bits_taken; // @[RocketTile.scala 130:32]
  assign frontend_io_cpu_bht_update_bits_mispredict = core_io_imem_bht_update_bits_mispredict; // @[RocketTile.scala 130:32]
  assign frontend_io_cpu_flush_icache = core_io_imem_flush_icache; // @[RocketTile.scala 130:32]
  assign frontend_io_ptw_req_ready = ptw_io_requestor_1_req_ready; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_resp_valid = ptw_io_requestor_1_resp_valid; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_resp_bits_ae = ptw_io_requestor_1_resp_bits_ae; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_resp_bits_pte_ppn = ptw_io_requestor_1_resp_bits_pte_ppn; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_resp_bits_pte_d = ptw_io_requestor_1_resp_bits_pte_d; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_resp_bits_pte_a = ptw_io_requestor_1_resp_bits_pte_a; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_resp_bits_pte_g = ptw_io_requestor_1_resp_bits_pte_g; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_resp_bits_pte_u = ptw_io_requestor_1_resp_bits_pte_u; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_resp_bits_pte_x = ptw_io_requestor_1_resp_bits_pte_x; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_resp_bits_pte_w = ptw_io_requestor_1_resp_bits_pte_w; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_resp_bits_pte_r = ptw_io_requestor_1_resp_bits_pte_r; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_resp_bits_pte_v = ptw_io_requestor_1_resp_bits_pte_v; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_resp_bits_level = ptw_io_requestor_1_resp_bits_level; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_resp_bits_homogeneous = ptw_io_requestor_1_resp_bits_homogeneous; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_ptbr_mode = ptw_io_requestor_1_ptbr_mode; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_status_prv = ptw_io_requestor_1_status_prv; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_0_cfg_l = ptw_io_requestor_1_pmp_0_cfg_l; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_0_cfg_a = ptw_io_requestor_1_pmp_0_cfg_a; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_0_cfg_x = ptw_io_requestor_1_pmp_0_cfg_x; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_0_cfg_w = ptw_io_requestor_1_pmp_0_cfg_w; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_0_cfg_r = ptw_io_requestor_1_pmp_0_cfg_r; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_0_addr = ptw_io_requestor_1_pmp_0_addr; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_0_mask = ptw_io_requestor_1_pmp_0_mask; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_1_cfg_l = ptw_io_requestor_1_pmp_1_cfg_l; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_1_cfg_a = ptw_io_requestor_1_pmp_1_cfg_a; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_1_cfg_x = ptw_io_requestor_1_pmp_1_cfg_x; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_1_cfg_w = ptw_io_requestor_1_pmp_1_cfg_w; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_1_cfg_r = ptw_io_requestor_1_pmp_1_cfg_r; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_1_addr = ptw_io_requestor_1_pmp_1_addr; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_1_mask = ptw_io_requestor_1_pmp_1_mask; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_2_cfg_l = ptw_io_requestor_1_pmp_2_cfg_l; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_2_cfg_a = ptw_io_requestor_1_pmp_2_cfg_a; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_2_cfg_x = ptw_io_requestor_1_pmp_2_cfg_x; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_2_cfg_w = ptw_io_requestor_1_pmp_2_cfg_w; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_2_cfg_r = ptw_io_requestor_1_pmp_2_cfg_r; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_2_addr = ptw_io_requestor_1_pmp_2_addr; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_2_mask = ptw_io_requestor_1_pmp_2_mask; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_3_cfg_l = ptw_io_requestor_1_pmp_3_cfg_l; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_3_cfg_a = ptw_io_requestor_1_pmp_3_cfg_a; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_3_cfg_x = ptw_io_requestor_1_pmp_3_cfg_x; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_3_cfg_w = ptw_io_requestor_1_pmp_3_cfg_w; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_3_cfg_r = ptw_io_requestor_1_pmp_3_cfg_r; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_3_addr = ptw_io_requestor_1_pmp_3_addr; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_3_mask = ptw_io_requestor_1_pmp_3_mask; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_4_cfg_l = ptw_io_requestor_1_pmp_4_cfg_l; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_4_cfg_a = ptw_io_requestor_1_pmp_4_cfg_a; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_4_cfg_x = ptw_io_requestor_1_pmp_4_cfg_x; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_4_cfg_w = ptw_io_requestor_1_pmp_4_cfg_w; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_4_cfg_r = ptw_io_requestor_1_pmp_4_cfg_r; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_4_addr = ptw_io_requestor_1_pmp_4_addr; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_4_mask = ptw_io_requestor_1_pmp_4_mask; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_5_cfg_l = ptw_io_requestor_1_pmp_5_cfg_l; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_5_cfg_a = ptw_io_requestor_1_pmp_5_cfg_a; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_5_cfg_x = ptw_io_requestor_1_pmp_5_cfg_x; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_5_cfg_w = ptw_io_requestor_1_pmp_5_cfg_w; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_5_cfg_r = ptw_io_requestor_1_pmp_5_cfg_r; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_5_addr = ptw_io_requestor_1_pmp_5_addr; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_5_mask = ptw_io_requestor_1_pmp_5_mask; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_6_cfg_l = ptw_io_requestor_1_pmp_6_cfg_l; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_6_cfg_a = ptw_io_requestor_1_pmp_6_cfg_a; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_6_cfg_x = ptw_io_requestor_1_pmp_6_cfg_x; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_6_cfg_w = ptw_io_requestor_1_pmp_6_cfg_w; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_6_cfg_r = ptw_io_requestor_1_pmp_6_cfg_r; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_6_addr = ptw_io_requestor_1_pmp_6_addr; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_6_mask = ptw_io_requestor_1_pmp_6_mask; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_7_cfg_l = ptw_io_requestor_1_pmp_7_cfg_l; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_7_cfg_a = ptw_io_requestor_1_pmp_7_cfg_a; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_7_cfg_x = ptw_io_requestor_1_pmp_7_cfg_x; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_7_cfg_w = ptw_io_requestor_1_pmp_7_cfg_w; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_7_cfg_r = ptw_io_requestor_1_pmp_7_cfg_r; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_7_addr = ptw_io_requestor_1_pmp_7_addr; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_pmp_7_mask = ptw_io_requestor_1_pmp_7_mask; // @[RocketTile.scala 169:20]
  assign frontend_io_ptw_vpoffset_bits_value = ptw_io_requestor_1_vpoffset_bits_value; // @[RocketTile.scala 169:20]
  assign buffer_clock = clock;
  assign buffer_reset = reset;
  assign buffer_auto_in_a_valid = tlMasterXbar_auto_out_a_valid; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_a_bits_opcode = tlMasterXbar_auto_out_a_bits_opcode; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_a_bits_param = tlMasterXbar_auto_out_a_bits_param; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_a_bits_size = tlMasterXbar_auto_out_a_bits_size; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_a_bits_source = tlMasterXbar_auto_out_a_bits_source; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_a_bits_address = tlMasterXbar_auto_out_a_bits_address; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_a_bits_mask = tlMasterXbar_auto_out_a_bits_mask; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_a_bits_data = tlMasterXbar_auto_out_a_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_a_bits_corrupt = tlMasterXbar_auto_out_a_bits_corrupt; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_b_ready = tlMasterXbar_auto_out_b_ready; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_c_valid = tlMasterXbar_auto_out_c_valid; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_c_bits_opcode = tlMasterXbar_auto_out_c_bits_opcode; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_c_bits_param = tlMasterXbar_auto_out_c_bits_param; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_c_bits_size = tlMasterXbar_auto_out_c_bits_size; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_c_bits_source = tlMasterXbar_auto_out_c_bits_source; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_c_bits_address = tlMasterXbar_auto_out_c_bits_address; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_c_bits_data = tlMasterXbar_auto_out_c_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_d_ready = tlMasterXbar_auto_out_d_ready; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_e_valid = tlMasterXbar_auto_out_e_valid; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_e_bits_sink = tlMasterXbar_auto_out_e_bits_sink; // @[LazyModule.scala 167:57]
  assign buffer_auto_out_a_ready = auto_tl_master_xing_out_a_ready; // @[LazyModule.scala 167:31]
  assign buffer_auto_out_b_valid = auto_tl_master_xing_out_b_valid; // @[LazyModule.scala 167:31]
  assign buffer_auto_out_b_bits_opcode = auto_tl_master_xing_out_b_bits_opcode; // @[LazyModule.scala 167:31]
  assign buffer_auto_out_b_bits_param = auto_tl_master_xing_out_b_bits_param; // @[LazyModule.scala 167:31]
  assign buffer_auto_out_b_bits_size = auto_tl_master_xing_out_b_bits_size; // @[LazyModule.scala 167:31]
  assign buffer_auto_out_b_bits_source = auto_tl_master_xing_out_b_bits_source; // @[LazyModule.scala 167:31]
  assign buffer_auto_out_b_bits_address = auto_tl_master_xing_out_b_bits_address; // @[LazyModule.scala 167:31]
  assign buffer_auto_out_b_bits_mask = auto_tl_master_xing_out_b_bits_mask; // @[LazyModule.scala 167:31]
  assign buffer_auto_out_b_bits_corrupt = auto_tl_master_xing_out_b_bits_corrupt; // @[LazyModule.scala 167:31]
  assign buffer_auto_out_c_ready = auto_tl_master_xing_out_c_ready; // @[LazyModule.scala 167:31]
  assign buffer_auto_out_d_valid = auto_tl_master_xing_out_d_valid; // @[LazyModule.scala 167:31]
  assign buffer_auto_out_d_bits_opcode = auto_tl_master_xing_out_d_bits_opcode; // @[LazyModule.scala 167:31]
  assign buffer_auto_out_d_bits_param = auto_tl_master_xing_out_d_bits_param; // @[LazyModule.scala 167:31]
  assign buffer_auto_out_d_bits_size = auto_tl_master_xing_out_d_bits_size; // @[LazyModule.scala 167:31]
  assign buffer_auto_out_d_bits_source = auto_tl_master_xing_out_d_bits_source; // @[LazyModule.scala 167:31]
  assign buffer_auto_out_d_bits_sink = auto_tl_master_xing_out_d_bits_sink; // @[LazyModule.scala 167:31]
  assign buffer_auto_out_d_bits_denied = auto_tl_master_xing_out_d_bits_denied; // @[LazyModule.scala 167:31]
  assign buffer_auto_out_d_bits_data = auto_tl_master_xing_out_d_bits_data; // @[LazyModule.scala 167:31]
  assign buffer_auto_out_d_bits_corrupt = auto_tl_master_xing_out_d_bits_corrupt; // @[LazyModule.scala 167:31]
  assign buffer_auto_out_e_ready = auto_tl_master_xing_out_e_ready; // @[LazyModule.scala 167:31]
  assign intsink_clock = clock;
  assign intsink_auto_in_sync_0 = auto_intsink_in_sync_0; // @[LazyModule.scala 173:31]
  assign intsink_1_auto_in_sync_0 = auto_int_in_xing_in_0_sync_0; // @[LazyModule.scala 167:57]
  assign intsink_1_auto_in_sync_1 = auto_int_in_xing_in_0_sync_1; // @[LazyModule.scala 167:57]
  assign intsink_2_auto_in_sync_0 = auto_int_in_xing_in_1_sync_0; // @[LazyModule.scala 167:57]
  assign intsink_3_auto_in_sync_0 = auto_int_in_xing_in_2_sync_0; // @[LazyModule.scala 167:57]
  assign fpuOpt_clock = clock;
  assign fpuOpt_reset = reset;
  assign fpuOpt_io_inst = core_io_fpu_inst; // @[RocketTile.scala 135:39]
  assign fpuOpt_io_fromint_data = core_io_fpu_fromint_data; // @[RocketTile.scala 135:39]
  assign fpuOpt_io_fcsr_rm = core_io_fpu_fcsr_rm; // @[RocketTile.scala 135:39]
  assign fpuOpt_io_dmem_resp_val = core_io_fpu_dmem_resp_val; // @[RocketTile.scala 135:39]
  assign fpuOpt_io_dmem_resp_type = core_io_fpu_dmem_resp_type; // @[RocketTile.scala 135:39]
  assign fpuOpt_io_dmem_resp_tag = core_io_fpu_dmem_resp_tag; // @[RocketTile.scala 135:39]
  assign fpuOpt_io_dmem_resp_data = core_io_fpu_dmem_resp_data; // @[RocketTile.scala 135:39]
  assign fpuOpt_io_valid = core_io_fpu_valid; // @[RocketTile.scala 135:39]
  assign fpuOpt_io_killx = core_io_fpu_killx; // @[RocketTile.scala 135:39]
  assign fpuOpt_io_killm = core_io_fpu_killm; // @[RocketTile.scala 135:39]
  assign dcacheArb_clock = clock;
  assign dcacheArb_io_requestor_0_req_valid = ptw_io_mem_req_valid; // @[RocketTile.scala 168:26]
  assign dcacheArb_io_requestor_0_req_bits_addr = ptw_io_mem_req_bits_addr; // @[RocketTile.scala 168:26]
  assign dcacheArb_io_requestor_0_s1_kill = ptw_io_mem_s1_kill; // @[RocketTile.scala 168:26]
  assign dcacheArb_io_requestor_1_req_valid = core_io_dmem_req_valid; // @[RocketTile.scala 168:26]
  assign dcacheArb_io_requestor_1_req_bits_addr = core_io_dmem_req_bits_addr; // @[RocketTile.scala 168:26]
  assign dcacheArb_io_requestor_1_req_bits_tag = core_io_dmem_req_bits_tag; // @[RocketTile.scala 168:26]
  assign dcacheArb_io_requestor_1_req_bits_cmd = core_io_dmem_req_bits_cmd; // @[RocketTile.scala 168:26]
  assign dcacheArb_io_requestor_1_req_bits_typ = core_io_dmem_req_bits_typ; // @[RocketTile.scala 168:26]
  assign dcacheArb_io_requestor_1_s1_kill = core_io_dmem_s1_kill; // @[RocketTile.scala 168:26]
  assign dcacheArb_io_requestor_1_s1_data_data = core_io_dmem_s1_data_data; // @[RocketTile.scala 168:26]
  assign dcacheArb_io_requestor_1_keep_clock_enabled = core_io_dmem_keep_clock_enabled; // @[RocketTile.scala 168:26]
  assign dcacheArb_io_mem_req_ready = dcache_io_cpu_req_ready; // @[HellaCache.scala 228:30]
  assign dcacheArb_io_mem_s2_nack = dcache_io_cpu_s2_nack; // @[HellaCache.scala 228:30]
  assign dcacheArb_io_mem_resp_valid = dcache_io_cpu_resp_valid; // @[HellaCache.scala 228:30]
  assign dcacheArb_io_mem_resp_bits_tag = dcache_io_cpu_resp_bits_tag; // @[HellaCache.scala 228:30]
  assign dcacheArb_io_mem_resp_bits_typ = dcache_io_cpu_resp_bits_typ; // @[HellaCache.scala 228:30]
  assign dcacheArb_io_mem_resp_bits_data = dcache_io_cpu_resp_bits_data; // @[HellaCache.scala 228:30]
  assign dcacheArb_io_mem_resp_bits_replay = dcache_io_cpu_resp_bits_replay; // @[HellaCache.scala 228:30]
  assign dcacheArb_io_mem_resp_bits_has_data = dcache_io_cpu_resp_bits_has_data; // @[HellaCache.scala 228:30]
  assign dcacheArb_io_mem_resp_bits_data_word_bypass = dcache_io_cpu_resp_bits_data_word_bypass; // @[HellaCache.scala 228:30]
  assign dcacheArb_io_mem_replay_next = dcache_io_cpu_replay_next; // @[HellaCache.scala 228:30]
  assign dcacheArb_io_mem_s2_xcpt_ma_ld = dcache_io_cpu_s2_xcpt_ma_ld; // @[HellaCache.scala 228:30]
  assign dcacheArb_io_mem_s2_xcpt_ma_st = dcache_io_cpu_s2_xcpt_ma_st; // @[HellaCache.scala 228:30]
  assign dcacheArb_io_mem_s2_xcpt_pf_ld = dcache_io_cpu_s2_xcpt_pf_ld; // @[HellaCache.scala 228:30]
  assign dcacheArb_io_mem_s2_xcpt_pf_st = dcache_io_cpu_s2_xcpt_pf_st; // @[HellaCache.scala 228:30]
  assign dcacheArb_io_mem_s2_xcpt_ae_ld = dcache_io_cpu_s2_xcpt_ae_ld; // @[HellaCache.scala 228:30]
  assign dcacheArb_io_mem_s2_xcpt_ae_st = dcache_io_cpu_s2_xcpt_ae_st; // @[HellaCache.scala 228:30]
  assign dcacheArb_io_mem_ordered = dcache_io_cpu_ordered; // @[HellaCache.scala 228:30]
  assign dcacheArb_io_mem_perf_grant = dcache_io_cpu_perf_grant; // @[HellaCache.scala 228:30]
  assign dcacheArb_io_mem_clock_enabled = dcache_io_cpu_clock_enabled; // @[HellaCache.scala 228:30]
  assign ptw_clock = clock;
  assign ptw_reset = reset;
  assign ptw_io_requestor_0_req_valid = dcache_io_ptw_req_valid; // @[RocketTile.scala 169:20]
  assign ptw_io_requestor_0_req_bits_bits_addr = dcache_io_ptw_req_bits_bits_addr; // @[RocketTile.scala 169:20]
  assign ptw_io_requestor_1_req_valid = frontend_io_ptw_req_valid; // @[RocketTile.scala 169:20]
  assign ptw_io_requestor_1_req_bits_valid = frontend_io_ptw_req_bits_valid; // @[RocketTile.scala 169:20]
  assign ptw_io_requestor_1_req_bits_bits_addr = frontend_io_ptw_req_bits_bits_addr; // @[RocketTile.scala 169:20]
  assign ptw_io_mem_req_ready = dcacheArb_io_requestor_0_req_ready; // @[RocketTile.scala 168:26]
  assign ptw_io_mem_s2_nack = dcacheArb_io_requestor_0_s2_nack; // @[RocketTile.scala 168:26]
  assign ptw_io_mem_resp_valid = dcacheArb_io_requestor_0_resp_valid; // @[RocketTile.scala 168:26]
  assign ptw_io_mem_resp_bits_data_word_bypass = dcacheArb_io_requestor_0_resp_bits_data_word_bypass; // @[RocketTile.scala 168:26]
  assign ptw_io_mem_s2_xcpt_ae_ld = dcacheArb_io_requestor_0_s2_xcpt_ae_ld; // @[RocketTile.scala 168:26]
  assign ptw_io_dpath_ptbr_mode = core_io_ptw_ptbr_mode; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_ptbr_ppn = core_io_ptw_ptbr_ppn; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_sfence_valid = core_io_ptw_sfence_valid; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_sfence_bits_rs1 = core_io_ptw_sfence_bits_rs1; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_status_dprv = core_io_ptw_status_dprv; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_status_prv = core_io_ptw_status_prv; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_status_mxr = core_io_ptw_status_mxr; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_status_sum = core_io_ptw_status_sum; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_0_cfg_l = core_io_ptw_pmp_0_cfg_l; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_0_cfg_a = core_io_ptw_pmp_0_cfg_a; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_0_cfg_x = core_io_ptw_pmp_0_cfg_x; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_0_cfg_w = core_io_ptw_pmp_0_cfg_w; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_0_cfg_r = core_io_ptw_pmp_0_cfg_r; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_0_addr = core_io_ptw_pmp_0_addr; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_0_mask = core_io_ptw_pmp_0_mask; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_1_cfg_l = core_io_ptw_pmp_1_cfg_l; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_1_cfg_a = core_io_ptw_pmp_1_cfg_a; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_1_cfg_x = core_io_ptw_pmp_1_cfg_x; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_1_cfg_w = core_io_ptw_pmp_1_cfg_w; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_1_cfg_r = core_io_ptw_pmp_1_cfg_r; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_1_addr = core_io_ptw_pmp_1_addr; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_1_mask = core_io_ptw_pmp_1_mask; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_2_cfg_l = core_io_ptw_pmp_2_cfg_l; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_2_cfg_a = core_io_ptw_pmp_2_cfg_a; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_2_cfg_x = core_io_ptw_pmp_2_cfg_x; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_2_cfg_w = core_io_ptw_pmp_2_cfg_w; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_2_cfg_r = core_io_ptw_pmp_2_cfg_r; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_2_addr = core_io_ptw_pmp_2_addr; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_2_mask = core_io_ptw_pmp_2_mask; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_3_cfg_l = core_io_ptw_pmp_3_cfg_l; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_3_cfg_a = core_io_ptw_pmp_3_cfg_a; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_3_cfg_x = core_io_ptw_pmp_3_cfg_x; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_3_cfg_w = core_io_ptw_pmp_3_cfg_w; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_3_cfg_r = core_io_ptw_pmp_3_cfg_r; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_3_addr = core_io_ptw_pmp_3_addr; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_3_mask = core_io_ptw_pmp_3_mask; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_4_cfg_l = core_io_ptw_pmp_4_cfg_l; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_4_cfg_a = core_io_ptw_pmp_4_cfg_a; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_4_cfg_x = core_io_ptw_pmp_4_cfg_x; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_4_cfg_w = core_io_ptw_pmp_4_cfg_w; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_4_cfg_r = core_io_ptw_pmp_4_cfg_r; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_4_addr = core_io_ptw_pmp_4_addr; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_4_mask = core_io_ptw_pmp_4_mask; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_5_cfg_l = core_io_ptw_pmp_5_cfg_l; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_5_cfg_a = core_io_ptw_pmp_5_cfg_a; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_5_cfg_x = core_io_ptw_pmp_5_cfg_x; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_5_cfg_w = core_io_ptw_pmp_5_cfg_w; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_5_cfg_r = core_io_ptw_pmp_5_cfg_r; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_5_addr = core_io_ptw_pmp_5_addr; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_5_mask = core_io_ptw_pmp_5_mask; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_6_cfg_l = core_io_ptw_pmp_6_cfg_l; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_6_cfg_a = core_io_ptw_pmp_6_cfg_a; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_6_cfg_x = core_io_ptw_pmp_6_cfg_x; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_6_cfg_w = core_io_ptw_pmp_6_cfg_w; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_6_cfg_r = core_io_ptw_pmp_6_cfg_r; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_6_addr = core_io_ptw_pmp_6_addr; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_6_mask = core_io_ptw_pmp_6_mask; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_7_cfg_l = core_io_ptw_pmp_7_cfg_l; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_7_cfg_a = core_io_ptw_pmp_7_cfg_a; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_7_cfg_x = core_io_ptw_pmp_7_cfg_x; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_7_cfg_w = core_io_ptw_pmp_7_cfg_w; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_7_cfg_r = core_io_ptw_pmp_7_cfg_r; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_7_addr = core_io_ptw_pmp_7_addr; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pmp_7_mask = core_io_ptw_pmp_7_mask; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pcode_req_valid = core_io_ptw_pcode_req_valid; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pcode_req_bits_id = core_io_ptw_pcode_req_bits_id; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pcode_req_bits_value_base = core_io_ptw_pcode_req_bits_value_base; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pcode_req_bits_value_mask = core_io_ptw_pcode_req_bits_value_mask; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pcode_req_bits_value_valid = core_io_ptw_pcode_req_bits_value_valid; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_pcode_req_bits_value_locked = core_io_ptw_pcode_req_bits_value_locked; // @[RocketTile.scala 141:15]
  assign ptw_io_dpath_vpoffset_req_bits_value = core_io_ptw_vpoffset_req_bits_value; // @[RocketTile.scala 141:15]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_hartid = constants_hartid; // @[RocketTile.scala 127:18]
  assign core_io_interrupts_debug = intXbar_auto_int_out_0; // @[Interrupts.scala 75:93]
  assign core_io_interrupts_mtip = intXbar_auto_int_out_2; // @[Interrupts.scala 75:93]
  assign core_io_interrupts_msip = intXbar_auto_int_out_1; // @[Interrupts.scala 75:93]
  assign core_io_interrupts_meip = intXbar_auto_int_out_3; // @[Interrupts.scala 75:93]
  assign core_io_interrupts_seip = intXbar_auto_int_out_4; // @[Interrupts.scala 75:93]
  assign core_io_imem_resp_valid = frontend_io_cpu_resp_valid; // @[RocketTile.scala 130:32]
  assign core_io_imem_resp_bits_btb_taken = frontend_io_cpu_resp_bits_btb_taken; // @[RocketTile.scala 130:32]
  assign core_io_imem_resp_bits_btb_bridx = frontend_io_cpu_resp_bits_btb_bridx; // @[RocketTile.scala 130:32]
  assign core_io_imem_resp_bits_btb_entry = frontend_io_cpu_resp_bits_btb_entry; // @[RocketTile.scala 130:32]
  assign core_io_imem_resp_bits_btb_bht_history = frontend_io_cpu_resp_bits_btb_bht_history; // @[RocketTile.scala 130:32]
  assign core_io_imem_resp_bits_pc = frontend_io_cpu_resp_bits_pc; // @[RocketTile.scala 130:32]
  assign core_io_imem_resp_bits_data = frontend_io_cpu_resp_bits_data; // @[RocketTile.scala 130:32]
  assign core_io_imem_resp_bits_xcpt_pf_inst = frontend_io_cpu_resp_bits_xcpt_pf_inst; // @[RocketTile.scala 130:32]
  assign core_io_imem_resp_bits_xcpt_ae_inst = frontend_io_cpu_resp_bits_xcpt_ae_inst; // @[RocketTile.scala 130:32]
  assign core_io_imem_resp_bits_replay = frontend_io_cpu_resp_bits_replay; // @[RocketTile.scala 130:32]
  assign core_io_dmem_req_ready = dcacheArb_io_requestor_1_req_ready; // @[RocketTile.scala 168:26]
  assign core_io_dmem_s2_nack = dcacheArb_io_requestor_1_s2_nack; // @[RocketTile.scala 168:26]
  assign core_io_dmem_resp_valid = dcacheArb_io_requestor_1_resp_valid; // @[RocketTile.scala 168:26]
  assign core_io_dmem_resp_bits_tag = dcacheArb_io_requestor_1_resp_bits_tag; // @[RocketTile.scala 168:26]
  assign core_io_dmem_resp_bits_typ = dcacheArb_io_requestor_1_resp_bits_typ; // @[RocketTile.scala 168:26]
  assign core_io_dmem_resp_bits_data = dcacheArb_io_requestor_1_resp_bits_data; // @[RocketTile.scala 168:26]
  assign core_io_dmem_resp_bits_replay = dcacheArb_io_requestor_1_resp_bits_replay; // @[RocketTile.scala 168:26]
  assign core_io_dmem_resp_bits_has_data = dcacheArb_io_requestor_1_resp_bits_has_data; // @[RocketTile.scala 168:26]
  assign core_io_dmem_resp_bits_data_word_bypass = dcacheArb_io_requestor_1_resp_bits_data_word_bypass; // @[RocketTile.scala 168:26]
  assign core_io_dmem_replay_next = dcacheArb_io_requestor_1_replay_next; // @[RocketTile.scala 168:26]
  assign core_io_dmem_s2_xcpt_ma_ld = dcacheArb_io_requestor_1_s2_xcpt_ma_ld; // @[RocketTile.scala 168:26]
  assign core_io_dmem_s2_xcpt_ma_st = dcacheArb_io_requestor_1_s2_xcpt_ma_st; // @[RocketTile.scala 168:26]
  assign core_io_dmem_s2_xcpt_pf_ld = dcacheArb_io_requestor_1_s2_xcpt_pf_ld; // @[RocketTile.scala 168:26]
  assign core_io_dmem_s2_xcpt_pf_st = dcacheArb_io_requestor_1_s2_xcpt_pf_st; // @[RocketTile.scala 168:26]
  assign core_io_dmem_s2_xcpt_ae_ld = dcacheArb_io_requestor_1_s2_xcpt_ae_ld; // @[RocketTile.scala 168:26]
  assign core_io_dmem_s2_xcpt_ae_st = dcacheArb_io_requestor_1_s2_xcpt_ae_st; // @[RocketTile.scala 168:26]
  assign core_io_dmem_ordered = dcacheArb_io_requestor_1_ordered; // @[RocketTile.scala 168:26]
  assign core_io_dmem_perf_grant = dcacheArb_io_requestor_1_perf_grant; // @[RocketTile.scala 168:26]
  assign core_io_dmem_clock_enabled = dcacheArb_io_requestor_1_clock_enabled; // @[RocketTile.scala 168:26]
  assign core_io_fpu_fcsr_flags_valid = fpuOpt_io_fcsr_flags_valid; // @[RocketTile.scala 135:39]
  assign core_io_fpu_fcsr_flags_bits = fpuOpt_io_fcsr_flags_bits; // @[RocketTile.scala 135:39]
  assign core_io_fpu_store_data = fpuOpt_io_store_data; // @[RocketTile.scala 135:39]
  assign core_io_fpu_toint_data = fpuOpt_io_toint_data; // @[RocketTile.scala 135:39]
  assign core_io_fpu_fcsr_rdy = fpuOpt_io_fcsr_rdy; // @[RocketTile.scala 135:39]
  assign core_io_fpu_nack_mem = fpuOpt_io_nack_mem; // @[RocketTile.scala 135:39]
  assign core_io_fpu_illegal_rm = fpuOpt_io_illegal_rm; // @[RocketTile.scala 135:39]
  assign core_io_fpu_dec_wen = fpuOpt_io_dec_wen; // @[RocketTile.scala 135:39]
  assign core_io_fpu_dec_ren1 = fpuOpt_io_dec_ren1; // @[RocketTile.scala 135:39]
  assign core_io_fpu_dec_ren2 = fpuOpt_io_dec_ren2; // @[RocketTile.scala 135:39]
  assign core_io_fpu_dec_ren3 = fpuOpt_io_dec_ren3; // @[RocketTile.scala 135:39]
  assign core_io_fpu_sboard_set = fpuOpt_io_sboard_set; // @[RocketTile.scala 135:39]
  assign core_io_fpu_sboard_clr = fpuOpt_io_sboard_clr; // @[RocketTile.scala 135:39]
  assign core_io_fpu_sboard_clra = fpuOpt_io_sboard_clra; // @[RocketTile.scala 135:39]
  assign RocketTile_covSum = 30'h0;
  assign intsink_1_sum = RocketTile_covSum + intsink_1_io_covSum;
  assign intsink_sum = intsink_1_sum + intsink_io_covSum;
  assign dcache_sum = intsink_sum + dcache_io_covSum;
  assign dcacheArb_sum = dcache_sum + dcacheArb_io_covSum;
  assign intsink_2_sum = dcacheArb_sum + intsink_2_io_covSum;
  assign frontend_sum = intsink_2_sum + frontend_io_covSum;
  assign buffer_sum = frontend_sum + buffer_io_covSum;
  assign core_sum = buffer_sum + core_io_covSum;
  assign intsink_3_sum = core_sum + intsink_3_io_covSum;
  assign ptw_sum = intsink_3_sum + ptw_io_covSum;
  assign tlMasterXbar_sum = ptw_sum + tlMasterXbar_io_covSum;
  assign fpuOpt_sum = tlMasterXbar_sum + fpuOpt_io_covSum;
  assign intXbar_sum = fpuOpt_sum + intXbar_io_covSum;
  assign io_covSum = intXbar_sum;
  assign ptw_metaAssert_wire = ptw_metaAssert;
  assign intsink_1_metaAssert_wire = intsink_1_metaAssert;
  assign intsink_3_metaAssert_wire = intsink_3_metaAssert;
  assign intsink_metaAssert_wire = intsink_metaAssert;
  assign intXbar_metaAssert_wire = intXbar_metaAssert;
  assign tlMasterXbar_metaAssert_wire = tlMasterXbar_metaAssert;
  assign dcacheArb_metaAssert_wire = dcacheArb_metaAssert;
  assign frontend_metaAssert_wire = frontend_metaAssert;
  assign buffer_metaAssert_wire = buffer_metaAssert;
  assign fpuOpt_metaAssert_wire = fpuOpt_metaAssert;
  assign intsink_2_metaAssert_wire = intsink_2_metaAssert;
  assign core_metaAssert_wire = core_metaAssert;
  assign dcache_metaAssert_wire = dcache_metaAssert;
  assign RocketTile_or8 = frontend_metaAssert_wire | dcache_metaAssert_wire;
  assign RocketTile_or3 = tlMasterXbar_metaAssert_wire | RocketTile_or8;
  assign RocketTile_or10 = intXbar_metaAssert_wire | ptw_metaAssert_wire;
  assign RocketTile_or4 = fpuOpt_metaAssert_wire | RocketTile_or10;
  assign RocketTile_or1 = RocketTile_or3 | RocketTile_or4;
  assign RocketTile_or12 = intsink_2_metaAssert_wire | intsink_3_metaAssert_wire;
  assign RocketTile_or5 = intsink_1_metaAssert_wire | RocketTile_or12;
  assign RocketTile_or13 = core_metaAssert_wire | dcacheArb_metaAssert_wire;
  assign RocketTile_or14 = intsink_metaAssert_wire | buffer_metaAssert_wire;
  assign RocketTile_or6 = RocketTile_or13 | RocketTile_or14;
  assign RocketTile_or2 = RocketTile_or5 | RocketTile_or6;
  assign RocketTile_or0 = RocketTile_or1 | RocketTile_or2;
  assign metaAssert = RocketTile_metaAssert;
  assign intsink_metaReset = metaReset | intsink_halt;
  assign dcache_metaReset = metaReset | dcache_halt;
  assign dcacheArb_metaReset = metaReset | dcacheArb_halt;
  assign frontend_metaReset = metaReset | frontend_halt;
  assign buffer_metaReset = metaReset | buffer_halt;
  assign core_metaReset = metaReset | core_halt;
  assign ptw_metaReset = metaReset | ptw_halt;
  assign tlMasterXbar_metaReset = metaReset | tlMasterXbar_halt;
  assign fpuOpt_metaReset = metaReset | fpuOpt_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  RocketTile_metaAssert = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      RocketTile_metaAssert <= 1'h0;
    end else begin
      RocketTile_metaAssert <= RocketTile_metaAssert | RocketTile_or0;
    end
  end
endmodule
module TLXbar_8(
  input         clock,
  input         reset,
  output        auto_in_1_a_ready,
  input         auto_in_1_a_valid,
  input  [31:0] auto_in_1_a_bits_address,
  output        auto_in_1_d_valid,
  output [2:0]  auto_in_1_d_bits_opcode,
  output [3:0]  auto_in_1_d_bits_size,
  output [63:0] auto_in_1_d_bits_data,
  output        auto_in_1_d_bits_corrupt,
  output        auto_in_0_a_ready,
  input         auto_in_0_a_valid,
  input  [2:0]  auto_in_0_a_bits_opcode,
  input  [2:0]  auto_in_0_a_bits_param,
  input  [3:0]  auto_in_0_a_bits_size,
  input         auto_in_0_a_bits_source,
  input  [31:0] auto_in_0_a_bits_address,
  input  [7:0]  auto_in_0_a_bits_mask,
  input  [63:0] auto_in_0_a_bits_data,
  input         auto_in_0_b_ready,
  output        auto_in_0_b_valid,
  output [1:0]  auto_in_0_b_bits_param,
  output [3:0]  auto_in_0_b_bits_size,
  output        auto_in_0_b_bits_source,
  output [31:0] auto_in_0_b_bits_address,
  output        auto_in_0_c_ready,
  input         auto_in_0_c_valid,
  input  [2:0]  auto_in_0_c_bits_opcode,
  input  [2:0]  auto_in_0_c_bits_param,
  input  [3:0]  auto_in_0_c_bits_size,
  input         auto_in_0_c_bits_source,
  input  [31:0] auto_in_0_c_bits_address,
  input  [63:0] auto_in_0_c_bits_data,
  input         auto_in_0_d_ready,
  output        auto_in_0_d_valid,
  output [2:0]  auto_in_0_d_bits_opcode,
  output [1:0]  auto_in_0_d_bits_param,
  output [3:0]  auto_in_0_d_bits_size,
  output        auto_in_0_d_bits_source,
  output [1:0]  auto_in_0_d_bits_sink,
  output        auto_in_0_d_bits_denied,
  output [63:0] auto_in_0_d_bits_data,
  output        auto_in_0_e_ready,
  input         auto_in_0_e_valid,
  input  [1:0]  auto_in_0_e_bits_sink,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [3:0]  auto_out_a_bits_size,
  output [1:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_a_bits_corrupt,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [2:0]  auto_out_b_bits_opcode,
  input  [1:0]  auto_out_b_bits_param,
  input  [3:0]  auto_out_b_bits_size,
  input  [1:0]  auto_out_b_bits_source,
  input  [31:0] auto_out_b_bits_address,
  input  [7:0]  auto_out_b_bits_mask,
  input         auto_out_b_bits_corrupt,
  input         auto_out_c_ready,
  output        auto_out_c_valid,
  output [2:0]  auto_out_c_bits_opcode,
  output [2:0]  auto_out_c_bits_param,
  output [3:0]  auto_out_c_bits_size,
  output [1:0]  auto_out_c_bits_source,
  output [31:0] auto_out_c_bits_address,
  output [63:0] auto_out_c_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_param,
  input  [3:0]  auto_out_d_bits_size,
  input  [1:0]  auto_out_d_bits_source,
  input  [1:0]  auto_out_d_bits_sink,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  input         auto_out_e_ready,
  output        auto_out_e_valid,
  output [1:0]  auto_out_e_bits_sink,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         TLMonitor_halt,
  input         TLMonitor_1_halt
);
  wire  TLMonitor_clock; // @[Nodes.scala 25:25]
  wire  TLMonitor_reset; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_a_ready; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_a_valid; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_a_bits_opcode; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_a_bits_param; // @[Nodes.scala 25:25]
  wire [3:0] TLMonitor_io_in_a_bits_size; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_a_bits_source; // @[Nodes.scala 25:25]
  wire [31:0] TLMonitor_io_in_a_bits_address; // @[Nodes.scala 25:25]
  wire [7:0] TLMonitor_io_in_a_bits_mask; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_b_ready; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_b_valid; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_b_bits_opcode; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_b_bits_param; // @[Nodes.scala 25:25]
  wire [3:0] TLMonitor_io_in_b_bits_size; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_b_bits_source; // @[Nodes.scala 25:25]
  wire [31:0] TLMonitor_io_in_b_bits_address; // @[Nodes.scala 25:25]
  wire [7:0] TLMonitor_io_in_b_bits_mask; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_b_bits_corrupt; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_c_ready; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_c_valid; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_c_bits_opcode; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_c_bits_param; // @[Nodes.scala 25:25]
  wire [3:0] TLMonitor_io_in_c_bits_size; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_c_bits_source; // @[Nodes.scala 25:25]
  wire [31:0] TLMonitor_io_in_c_bits_address; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_d_ready; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_d_valid; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_d_bits_opcode; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_d_bits_param; // @[Nodes.scala 25:25]
  wire [3:0] TLMonitor_io_in_d_bits_size; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_d_bits_source; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_d_bits_sink; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_d_bits_denied; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_d_bits_corrupt; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_e_ready; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_e_valid; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_e_bits_sink; // @[Nodes.scala 25:25]
  wire [29:0] TLMonitor_io_covSum; // @[Nodes.scala 25:25]
  wire  TLMonitor_metaAssert; // @[Nodes.scala 25:25]
  wire  TLMonitor_metaReset; // @[Nodes.scala 25:25]
  wire  TLMonitor_1_clock; // @[Nodes.scala 25:25]
  wire  TLMonitor_1_reset; // @[Nodes.scala 25:25]
  wire  TLMonitor_1_io_in_a_ready; // @[Nodes.scala 25:25]
  wire  TLMonitor_1_io_in_a_valid; // @[Nodes.scala 25:25]
  wire [31:0] TLMonitor_1_io_in_a_bits_address; // @[Nodes.scala 25:25]
  wire  TLMonitor_1_io_in_d_valid; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_1_io_in_d_bits_opcode; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_1_io_in_d_bits_param; // @[Nodes.scala 25:25]
  wire [3:0] TLMonitor_1_io_in_d_bits_size; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_1_io_in_d_bits_sink; // @[Nodes.scala 25:25]
  wire  TLMonitor_1_io_in_d_bits_denied; // @[Nodes.scala 25:25]
  wire  TLMonitor_1_io_in_d_bits_corrupt; // @[Nodes.scala 25:25]
  wire [29:0] TLMonitor_1_io_covSum; // @[Nodes.scala 25:25]
  wire  TLMonitor_1_metaAssert; // @[Nodes.scala 25:25]
  wire  TLMonitor_1_metaReset; // @[Nodes.scala 25:25]
  wire  requestBOI_0_0; // @[Parameters.scala 52:32]
  wire  requestDOI_0_0; // @[Parameters.scala 52:32]
  wire  requestDOI_0_1; // @[Parameters.scala 44:9]
  wire [26:0] _T_818; // @[package.scala 185:77]
  wire [8:0] _T_821; // @[Edges.scala 220:59]
  wire  _T_1001; // @[Mux.scala 19:72]
  reg [8:0] _T_1047; // @[Arbiter.scala 53:30]
  reg [31:0] _RAND_0;
  wire  _T_1048; // @[Arbiter.scala 54:28]
  wire  _T_1049; // @[Arbiter.scala 55:24]
  wire [1:0] _T_1050; // @[Cat.scala 30:58]
  wire  _T_1052; // @[Arbiter.scala 19:19]
  wire  _T_1054; // @[Arbiter.scala 19:12]
  reg [1:0] _T_1058; // @[Arbiter.scala 20:23]
  reg [31:0] _RAND_1;
  wire [1:0] _T_1060; // @[Arbiter.scala 21:28]
  wire [3:0] _T_1061; // @[Cat.scala 30:58]
  wire [3:0] _GEN_1; // @[package.scala 203:43]
  wire [3:0] _T_1063; // @[package.scala 203:43]
  wire [3:0] _T_1066; // @[Arbiter.scala 22:66]
  wire [3:0] _GEN_2; // @[Arbiter.scala 22:58]
  wire [3:0] _T_1067; // @[Arbiter.scala 22:58]
  wire [1:0] _T_1070; // @[Arbiter.scala 23:39]
  wire  _T_1072; // @[Arbiter.scala 24:27]
  wire  _T_1073; // @[Arbiter.scala 24:18]
  wire [1:0] _T_1074; // @[Arbiter.scala 25:29]
  wire [2:0] _T_1075; // @[package.scala 194:48]
  wire [1:0] _T_1077; // @[package.scala 194:43]
  wire  _T_1080; // @[Arbiter.scala 60:72]
  wire  _T_1081; // @[Arbiter.scala 60:72]
  wire  _T_1090; // @[Arbiter.scala 62:65]
  wire  _T_1091; // @[Arbiter.scala 62:65]
  wire  _T_1101; // @[Arbiter.scala 67:52]
  wire  _T_1107; // @[Arbiter.scala 68:59]
  wire  _T_1110; // @[Arbiter.scala 68:13]
  wire  _T_1112; // @[Arbiter.scala 70:31]
  wire  _T_1115; // @[Arbiter.scala 70:36]
  wire  _T_1117; // @[Arbiter.scala 70:14]
  reg  _T_1143_0; // @[Arbiter.scala 78:26]
  reg [31:0] _RAND_2;
  wire  _T_1174; // @[Mux.scala 19:72]
  reg  _T_1143_1; // @[Arbiter.scala 78:26]
  reg [31:0] _RAND_3;
  wire  _T_1175; // @[Mux.scala 19:72]
  wire  _T_1176; // @[Mux.scala 19:72]
  wire  out_0_a_valid; // @[Arbiter.scala 86:24]
  wire  _T_1122; // @[Decoupled.scala 37:37]
  wire [8:0] _GEN_3; // @[Arbiter.scala 75:52]
  wire [8:0] _T_1125; // @[Arbiter.scala 75:52]
  wire  _T_1154_0; // @[Arbiter.scala 79:25]
  wire  _T_1154_1; // @[Arbiter.scala 79:25]
  wire  _T_1162_0; // @[Arbiter.scala 82:24]
  wire  _T_1162_1; // @[Arbiter.scala 82:24]
  wire [1:0] in_0_a_bits_source; // @[Xbar.scala 109:18 Xbar.scala 114:17 Xbar.scala 115:29]
  wire [116:0] _T_1187; // @[Mux.scala 19:72]
  wire [116:0] _T_1188; // @[Mux.scala 19:72]
  wire [116:0] _T_1195; // @[Mux.scala 19:72]
  wire [116:0] _T_1196; // @[Mux.scala 19:72]
  wire [116:0] _T_1197; // @[Mux.scala 19:72]
  reg [2:0] TLXbar_8_state; // @[Register tracking TLXbar_8 state]
  reg [31:0] _RAND_4;
  reg  TLXbar_8_cov [0:7]; // @[Coverage map for TLXbar_8]
  reg [31:0] _RAND_5;
  wire  TLXbar_8_cov_read_data; // @[Coverage map for TLXbar_8]
  wire [2:0] TLXbar_8_cov_read_addr; // @[Coverage map for TLXbar_8]
  wire  TLXbar_8_cov_write_data; // @[Coverage map for TLXbar_8]
  wire [2:0] TLXbar_8_cov_write_addr; // @[Coverage map for TLXbar_8]
  wire  TLXbar_8_cov_write_mask; // @[Coverage map for TLXbar_8]
  wire  TLXbar_8_cov_write_en; // @[Coverage map for TLXbar_8]
  reg [29:0] TLXbar_8_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_6;
  wire [1:0] _T_1058_shl;
  wire [2:0] _T_1058_pad;
  wire [2:0] _T_1143_0_shl;
  wire [2:0] _T_1143_0_pad;
  wire [2:0] _T_1143_1_shl;
  wire [2:0] _T_1143_1_pad;
  wire [2:0] TLXbar_8_xor2;
  wire [2:0] TLXbar_8_xor0;
  wire [29:0] TLMonitor_sum;
  wire [29:0] TLMonitor_1_sum;
  wire  stopEn0;
  wire  stopEn1;
  wire  stopEn2;
  wire  TLMonitor_metaAssert_wire;
  wire  TLMonitor_1_metaAssert_wire;
  wire  TLXbar_8_or1;
  wire  TLXbar_8_or6;
  wire  TLXbar_8_or2;
  wire  TLXbar_8_or0;
  reg  TLXbar_8_metaAssert;
  reg [31:0] _RAND_7;
  TLMonitor_64 TLMonitor ( // @[Nodes.scala 25:25]
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_b_ready(TLMonitor_io_in_b_ready),
    .io_in_b_valid(TLMonitor_io_in_b_valid),
    .io_in_b_bits_opcode(TLMonitor_io_in_b_bits_opcode),
    .io_in_b_bits_param(TLMonitor_io_in_b_bits_param),
    .io_in_b_bits_size(TLMonitor_io_in_b_bits_size),
    .io_in_b_bits_source(TLMonitor_io_in_b_bits_source),
    .io_in_b_bits_address(TLMonitor_io_in_b_bits_address),
    .io_in_b_bits_mask(TLMonitor_io_in_b_bits_mask),
    .io_in_b_bits_corrupt(TLMonitor_io_in_b_bits_corrupt),
    .io_in_c_ready(TLMonitor_io_in_c_ready),
    .io_in_c_valid(TLMonitor_io_in_c_valid),
    .io_in_c_bits_opcode(TLMonitor_io_in_c_bits_opcode),
    .io_in_c_bits_param(TLMonitor_io_in_c_bits_param),
    .io_in_c_bits_size(TLMonitor_io_in_c_bits_size),
    .io_in_c_bits_source(TLMonitor_io_in_c_bits_source),
    .io_in_c_bits_address(TLMonitor_io_in_c_bits_address),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt),
    .io_in_e_ready(TLMonitor_io_in_e_ready),
    .io_in_e_valid(TLMonitor_io_in_e_valid),
    .io_in_e_bits_sink(TLMonitor_io_in_e_bits_sink),
    .io_covSum(TLMonitor_io_covSum),
    .metaAssert(TLMonitor_metaAssert),
    .metaReset(TLMonitor_metaReset)
  );
  TLMonitor_65 TLMonitor_1 ( // @[Nodes.scala 25:25]
    .clock(TLMonitor_1_clock),
    .reset(TLMonitor_1_reset),
    .io_in_a_ready(TLMonitor_1_io_in_a_ready),
    .io_in_a_valid(TLMonitor_1_io_in_a_valid),
    .io_in_a_bits_address(TLMonitor_1_io_in_a_bits_address),
    .io_in_d_valid(TLMonitor_1_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_1_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_1_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_1_io_in_d_bits_size),
    .io_in_d_bits_sink(TLMonitor_1_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_1_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_1_io_in_d_bits_corrupt),
    .io_covSum(TLMonitor_1_io_covSum),
    .metaAssert(TLMonitor_1_metaAssert),
    .metaReset(TLMonitor_1_metaReset)
  );
  assign requestBOI_0_0 = ~auto_out_b_bits_source[1]; // @[Parameters.scala 52:32]
  assign requestDOI_0_0 = ~auto_out_d_bits_source[1]; // @[Parameters.scala 52:32]
  assign requestDOI_0_1 = auto_out_d_bits_source == 2'h2; // @[Parameters.scala 44:9]
  assign _T_818 = 27'hfff << auto_in_0_a_bits_size; // @[package.scala 185:77]
  assign _T_821 = ~_T_818[11:3]; // @[Edges.scala 220:59]
  assign _T_1001 = requestDOI_0_0 & auto_in_0_d_ready; // @[Mux.scala 19:72]
  assign _T_1048 = _T_1047 == 9'h0; // @[Arbiter.scala 54:28]
  assign _T_1049 = _T_1048 & auto_out_a_ready; // @[Arbiter.scala 55:24]
  assign _T_1050 = {auto_in_1_a_valid,auto_in_0_a_valid}; // @[Cat.scala 30:58]
  assign _T_1052 = _T_1050 == _T_1050; // @[Arbiter.scala 19:19]
  assign _T_1054 = _T_1052 | reset; // @[Arbiter.scala 19:12]
  assign _T_1060 = _T_1050 & ~_T_1058; // @[Arbiter.scala 21:28]
  assign _T_1061 = {_T_1060,auto_in_1_a_valid,auto_in_0_a_valid}; // @[Cat.scala 30:58]
  assign _GEN_1 = {{1'd0}, _T_1061[3:1]}; // @[package.scala 203:43]
  assign _T_1063 = _T_1061 | _GEN_1; // @[package.scala 203:43]
  assign _T_1066 = {_T_1058, 2'h0}; // @[Arbiter.scala 22:66]
  assign _GEN_2 = {{1'd0}, _T_1063[3:1]}; // @[Arbiter.scala 22:58]
  assign _T_1067 = _GEN_2 | _T_1066; // @[Arbiter.scala 22:58]
  assign _T_1070 = _T_1067[3:2] & _T_1067[1:0]; // @[Arbiter.scala 23:39]
  assign _T_1072 = _T_1050 != 2'h0; // @[Arbiter.scala 24:27]
  assign _T_1073 = _T_1049 & _T_1072; // @[Arbiter.scala 24:18]
  assign _T_1074 = ~_T_1070 & _T_1050; // @[Arbiter.scala 25:29]
  assign _T_1075 = {_T_1074, 1'h0}; // @[package.scala 194:48]
  assign _T_1077 = _T_1074 | _T_1075[1:0]; // @[package.scala 194:43]
  assign _T_1080 = ~_T_1070[0]; // @[Arbiter.scala 60:72]
  assign _T_1081 = ~_T_1070[1]; // @[Arbiter.scala 60:72]
  assign _T_1090 = _T_1080 & auto_in_0_a_valid; // @[Arbiter.scala 62:65]
  assign _T_1091 = _T_1081 & auto_in_1_a_valid; // @[Arbiter.scala 62:65]
  assign _T_1101 = _T_1090 | _T_1091; // @[Arbiter.scala 67:52]
  assign _T_1107 = ~_T_1090 | ~_T_1091; // @[Arbiter.scala 68:59]
  assign _T_1110 = _T_1107 | reset; // @[Arbiter.scala 68:13]
  assign _T_1112 = auto_in_0_a_valid | auto_in_1_a_valid; // @[Arbiter.scala 70:31]
  assign _T_1115 = ~_T_1112 | _T_1101; // @[Arbiter.scala 70:36]
  assign _T_1117 = _T_1115 | reset; // @[Arbiter.scala 70:14]
  assign _T_1174 = _T_1143_0 & auto_in_0_a_valid; // @[Mux.scala 19:72]
  assign _T_1175 = _T_1143_1 & auto_in_1_a_valid; // @[Mux.scala 19:72]
  assign _T_1176 = _T_1174 | _T_1175; // @[Mux.scala 19:72]
  assign out_0_a_valid = _T_1048 ? _T_1112 : _T_1176; // @[Arbiter.scala 86:24]
  assign _T_1122 = auto_out_a_ready & out_0_a_valid; // @[Decoupled.scala 37:37]
  assign _GEN_3 = {{8'd0}, _T_1122}; // @[Arbiter.scala 75:52]
  assign _T_1125 = _T_1047 - _GEN_3; // @[Arbiter.scala 75:52]
  assign _T_1154_0 = _T_1048 ? _T_1090 : _T_1143_0; // @[Arbiter.scala 79:25]
  assign _T_1154_1 = _T_1048 ? _T_1091 : _T_1143_1; // @[Arbiter.scala 79:25]
  assign _T_1162_0 = _T_1048 ? _T_1080 : _T_1143_0; // @[Arbiter.scala 82:24]
  assign _T_1162_1 = _T_1048 ? _T_1081 : _T_1143_1; // @[Arbiter.scala 82:24]
  assign in_0_a_bits_source = {{1'd0}, auto_in_0_a_bits_source}; // @[Xbar.scala 109:18 Xbar.scala 114:17 Xbar.scala 115:29]
  assign _T_1187 = {auto_in_0_a_bits_opcode,auto_in_0_a_bits_param,auto_in_0_a_bits_size,in_0_a_bits_source,auto_in_0_a_bits_address,auto_in_0_a_bits_mask,auto_in_0_a_bits_data,1'h0}; // @[Mux.scala 19:72]
  assign _T_1188 = _T_1154_0 ? _T_1187 : 117'h0; // @[Mux.scala 19:72]
  assign _T_1195 = {12'h81a,auto_in_1_a_bits_address,8'hff,65'h0}; // @[Mux.scala 19:72]
  assign _T_1196 = _T_1154_1 ? _T_1195 : 117'h0; // @[Mux.scala 19:72]
  assign _T_1197 = _T_1188 | _T_1196; // @[Mux.scala 19:72]
  assign auto_in_1_a_ready = auto_out_a_ready & _T_1162_1; // @[LazyModule.scala 173:31]
  assign auto_in_1_d_valid = auto_out_d_valid & requestDOI_0_1; // @[LazyModule.scala 173:31]
  assign auto_in_1_d_bits_opcode = auto_out_d_bits_opcode; // @[LazyModule.scala 173:31]
  assign auto_in_1_d_bits_size = auto_out_d_bits_size; // @[LazyModule.scala 173:31]
  assign auto_in_1_d_bits_data = auto_out_d_bits_data; // @[LazyModule.scala 173:31]
  assign auto_in_1_d_bits_corrupt = auto_out_d_bits_corrupt; // @[LazyModule.scala 173:31]
  assign auto_in_0_a_ready = auto_out_a_ready & _T_1162_0; // @[LazyModule.scala 173:31]
  assign auto_in_0_b_valid = auto_out_b_valid & requestBOI_0_0; // @[LazyModule.scala 173:31]
  assign auto_in_0_b_bits_param = auto_out_b_bits_param; // @[LazyModule.scala 173:31]
  assign auto_in_0_b_bits_size = auto_out_b_bits_size; // @[LazyModule.scala 173:31]
  assign auto_in_0_b_bits_source = auto_out_b_bits_source[0]; // @[LazyModule.scala 173:31]
  assign auto_in_0_b_bits_address = auto_out_b_bits_address; // @[LazyModule.scala 173:31]
  assign auto_in_0_c_ready = auto_out_c_ready; // @[LazyModule.scala 173:31]
  assign auto_in_0_d_valid = auto_out_d_valid & requestDOI_0_0; // @[LazyModule.scala 173:31]
  assign auto_in_0_d_bits_opcode = auto_out_d_bits_opcode; // @[LazyModule.scala 173:31]
  assign auto_in_0_d_bits_param = auto_out_d_bits_param; // @[LazyModule.scala 173:31]
  assign auto_in_0_d_bits_size = auto_out_d_bits_size; // @[LazyModule.scala 173:31]
  assign auto_in_0_d_bits_source = auto_out_d_bits_source[0]; // @[LazyModule.scala 173:31]
  assign auto_in_0_d_bits_sink = auto_out_d_bits_sink; // @[LazyModule.scala 173:31]
  assign auto_in_0_d_bits_denied = auto_out_d_bits_denied; // @[LazyModule.scala 173:31]
  assign auto_in_0_d_bits_data = auto_out_d_bits_data; // @[LazyModule.scala 173:31]
  assign auto_in_0_e_ready = auto_out_e_ready; // @[LazyModule.scala 173:31]
  assign auto_out_a_valid = _T_1048 ? _T_1112 : _T_1176; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_opcode = _T_1197[116:114]; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_param = _T_1197[113:111]; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_size = _T_1197[110:107]; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_source = _T_1197[106:105]; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_address = _T_1197[104:73]; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_mask = _T_1197[72:65]; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_data = _T_1197[64:1]; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_corrupt = _T_1197[0]; // @[LazyModule.scala 173:49]
  assign auto_out_b_ready = requestBOI_0_0 & auto_in_0_b_ready; // @[LazyModule.scala 173:49]
  assign auto_out_c_valid = auto_in_0_c_valid; // @[LazyModule.scala 173:49]
  assign auto_out_c_bits_opcode = auto_in_0_c_bits_opcode; // @[LazyModule.scala 173:49]
  assign auto_out_c_bits_param = auto_in_0_c_bits_param; // @[LazyModule.scala 173:49]
  assign auto_out_c_bits_size = auto_in_0_c_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_c_bits_source = {{1'd0}, auto_in_0_c_bits_source}; // @[LazyModule.scala 173:49]
  assign auto_out_c_bits_address = auto_in_0_c_bits_address; // @[LazyModule.scala 173:49]
  assign auto_out_c_bits_data = auto_in_0_c_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_d_ready = _T_1001 | requestDOI_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_e_valid = auto_in_0_e_valid; // @[LazyModule.scala 173:49]
  assign auto_out_e_bits_sink = auto_in_0_e_bits_sink; // @[LazyModule.scala 173:49]
  assign TLMonitor_clock = clock;
  assign TLMonitor_reset = reset;
  assign TLMonitor_io_in_a_ready = auto_out_a_ready & _T_1162_0; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_valid = auto_in_0_a_valid; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_opcode = auto_in_0_a_bits_opcode; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_param = auto_in_0_a_bits_param; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_size = auto_in_0_a_bits_size; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_source = auto_in_0_a_bits_source; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_address = auto_in_0_a_bits_address; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_mask = auto_in_0_a_bits_mask; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_ready = auto_in_0_b_ready; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_valid = auto_out_b_valid & requestBOI_0_0; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_opcode = auto_out_b_bits_opcode; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_param = auto_out_b_bits_param; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_size = auto_out_b_bits_size; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_source = auto_out_b_bits_source[0]; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_address = auto_out_b_bits_address; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_mask = auto_out_b_bits_mask; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_corrupt = auto_out_b_bits_corrupt; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_ready = auto_out_c_ready; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_valid = auto_in_0_c_valid; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_bits_opcode = auto_in_0_c_bits_opcode; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_bits_param = auto_in_0_c_bits_param; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_bits_size = auto_in_0_c_bits_size; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_bits_source = auto_in_0_c_bits_source; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_bits_address = auto_in_0_c_bits_address; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_ready = auto_in_0_d_ready; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_valid = auto_out_d_valid & requestDOI_0_0; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_source = auto_out_d_bits_source[0]; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_e_ready = auto_out_e_ready; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_e_valid = auto_in_0_e_valid; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_e_bits_sink = auto_in_0_e_bits_sink; // @[Nodes.scala 26:19]
  assign TLMonitor_1_clock = clock;
  assign TLMonitor_1_reset = reset;
  assign TLMonitor_1_io_in_a_ready = auto_out_a_ready & _T_1162_1; // @[Nodes.scala 26:19]
  assign TLMonitor_1_io_in_a_valid = auto_in_1_a_valid; // @[Nodes.scala 26:19]
  assign TLMonitor_1_io_in_a_bits_address = auto_in_1_a_bits_address; // @[Nodes.scala 26:19]
  assign TLMonitor_1_io_in_d_valid = auto_out_d_valid & requestDOI_0_1; // @[Nodes.scala 26:19]
  assign TLMonitor_1_io_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 26:19]
  assign TLMonitor_1_io_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 26:19]
  assign TLMonitor_1_io_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 26:19]
  assign TLMonitor_1_io_in_d_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 26:19]
  assign TLMonitor_1_io_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 26:19]
  assign TLMonitor_1_io_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 26:19]
  assign TLXbar_8_cov_read_addr = TLXbar_8_state;
  assign TLXbar_8_cov_read_data = TLXbar_8_cov[TLXbar_8_cov_read_addr]; // @[Coverage map for TLXbar_8]
  assign TLXbar_8_cov_write_data = 1'h1;
  assign TLXbar_8_cov_write_addr = TLXbar_8_state;
  assign TLXbar_8_cov_write_mask = 1'h1;
  assign TLXbar_8_cov_write_en = 1'h1;
  assign _T_1058_shl = _T_1058;
  assign _T_1058_pad = {1'h0,_T_1058_shl};
  assign _T_1143_0_shl = {_T_1143_0, 2'h0};
  assign _T_1143_0_pad = _T_1143_0_shl;
  assign _T_1143_1_shl = {_T_1143_1, 2'h0};
  assign _T_1143_1_pad = _T_1143_1_shl;
  assign TLXbar_8_xor2 = _T_1143_0_pad ^ _T_1143_1_pad;
  assign TLXbar_8_xor0 = _T_1058_pad ^ TLXbar_8_xor2;
  assign TLMonitor_sum = TLXbar_8_covSum + TLMonitor_io_covSum;
  assign TLMonitor_1_sum = TLMonitor_sum + TLMonitor_1_io_covSum;
  assign io_covSum = TLMonitor_1_sum;
  assign stopEn0 = ~_T_1054;
  assign stopEn1 = ~_T_1110;
  assign stopEn2 = ~_T_1117;
  assign TLMonitor_metaAssert_wire = TLMonitor_metaAssert;
  assign TLMonitor_1_metaAssert_wire = TLMonitor_1_metaAssert;
  assign TLXbar_8_or1 = stopEn0 | stopEn1;
  assign TLXbar_8_or6 = TLMonitor_metaAssert_wire | TLMonitor_1_metaAssert_wire;
  assign TLXbar_8_or2 = stopEn2 | TLXbar_8_or6;
  assign TLXbar_8_or0 = TLXbar_8_or1 | TLXbar_8_or2;
  assign metaAssert = TLXbar_8_metaAssert;
  assign TLMonitor_metaReset = metaReset | TLMonitor_halt;
  assign TLMonitor_1_metaReset = metaReset | TLMonitor_1_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1047 = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1058 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1143_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1143_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  TLXbar_8_state = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    TLXbar_8_cov[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  TLXbar_8_covSum = _RAND_6[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  TLXbar_8_metaAssert = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      _T_1047 <= 9'h0;
    end else if (reset) begin
      _T_1047 <= 9'h0;
    end else if (_T_1049) begin
      if (_T_1090) begin
        if (~auto_in_0_a_bits_opcode[2]) begin
          _T_1047 <= _T_821;
        end else begin
          _T_1047 <= 9'h0;
        end
      end else begin
        _T_1047 <= 9'h0;
      end
    end else begin
      _T_1047 <= _T_1125;
    end
    if (metaReset) begin
      _T_1058 <= 2'h0;
    end else if (reset) begin
      _T_1058 <= 2'h3;
    end else if (_T_1073) begin
      _T_1058 <= _T_1077;
    end
    if (metaReset) begin
      _T_1143_0 <= 1'h0;
    end else if (reset) begin
      _T_1143_0 <= 1'h0;
    end else if (_T_1048) begin
      _T_1143_0 <= _T_1090;
    end
    if (metaReset) begin
      _T_1143_1 <= 1'h0;
    end else if (reset) begin
      _T_1143_1 <= 1'h0;
    end else if (_T_1048) begin
      _T_1143_1 <= _T_1091;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_1054) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n"); // @[Arbiter.scala 19:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_1054) begin
          $fatal; // @[Arbiter.scala 19:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_1110) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Arbiter.scala 68:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_1110) begin
          $fatal; // @[Arbiter.scala 68:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_1117) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:70 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n"); // @[Arbiter.scala 70:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_1117) begin
          $fatal; // @[Arbiter.scala 70:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    TLXbar_8_state <= TLXbar_8_xor0;
    if (!(TLXbar_8_cov_read_data)) begin
      TLXbar_8_covSum <= TLXbar_8_covSum + 1'h1;
    end
    if (metaReset) begin
      TLXbar_8_metaAssert <= 1'h0;
    end else begin
      TLXbar_8_metaAssert <= TLXbar_8_metaAssert | TLXbar_8_or0;
    end
  end
  always @(posedge clock) begin
    if(TLXbar_8_cov_write_en & TLXbar_8_cov_write_mask) begin
      TLXbar_8_cov[TLXbar_8_cov_write_addr] <= TLXbar_8_cov_write_data; // @[Coverage map for TLXbar_8]
    end
  end
endmodule
module IntXbar_1(
  input         auto_int_in_3_0,
  input         auto_int_in_2_0,
  input         auto_int_in_1_0,
  input         auto_int_in_1_1,
  input         auto_int_in_0_0,
  output        auto_int_out_0,
  output        auto_int_out_1,
  output        auto_int_out_2,
  output        auto_int_out_3,
  output        auto_int_out_4,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [29:0] IntXbar_1_covSum;
  assign auto_int_out_0 = auto_int_in_0_0; // @[LazyModule.scala 173:49]
  assign auto_int_out_1 = auto_int_in_1_0; // @[LazyModule.scala 173:49]
  assign auto_int_out_2 = auto_int_in_1_1; // @[LazyModule.scala 173:49]
  assign auto_int_out_3 = auto_int_in_2_0; // @[LazyModule.scala 173:49]
  assign auto_int_out_4 = auto_int_in_3_0; // @[LazyModule.scala 173:49]
  assign IntXbar_1_covSum = 30'h0;
  assign io_covSum = IntXbar_1_covSum;
  assign metaAssert = 1'h0;
endmodule
module DCache(
  input         gated_clock,
  input         reset,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [3:0]  auto_out_a_bits_size,
  output        auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [1:0]  auto_out_b_bits_param,
  input  [3:0]  auto_out_b_bits_size,
  input         auto_out_b_bits_source,
  input  [31:0] auto_out_b_bits_address,
  input         auto_out_c_ready,
  output        auto_out_c_valid,
  output [2:0]  auto_out_c_bits_opcode,
  output [2:0]  auto_out_c_bits_param,
  output [3:0]  auto_out_c_bits_size,
  output        auto_out_c_bits_source,
  output [31:0] auto_out_c_bits_address,
  output [63:0] auto_out_c_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_param,
  input  [3:0]  auto_out_d_bits_size,
  input         auto_out_d_bits_source,
  input  [1:0]  auto_out_d_bits_sink,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_e_ready,
  output        auto_out_e_valid,
  output [1:0]  auto_out_e_bits_sink,
  output        io_cpu_req_ready,
  input         io_cpu_req_valid,
  input  [39:0] io_cpu_req_bits_addr,
  input  [6:0]  io_cpu_req_bits_tag,
  input  [4:0]  io_cpu_req_bits_cmd,
  input  [2:0]  io_cpu_req_bits_typ,
  input         io_cpu_req_bits_phys,
  input         io_cpu_s1_kill,
  input  [63:0] io_cpu_s1_data_data,
  output        io_cpu_s2_nack,
  output        io_cpu_resp_valid,
  output [6:0]  io_cpu_resp_bits_tag,
  output [2:0]  io_cpu_resp_bits_typ,
  output [63:0] io_cpu_resp_bits_data,
  output        io_cpu_resp_bits_replay,
  output        io_cpu_resp_bits_has_data,
  output [63:0] io_cpu_resp_bits_data_word_bypass,
  output        io_cpu_replay_next,
  output        io_cpu_s2_xcpt_ma_ld,
  output        io_cpu_s2_xcpt_ma_st,
  output        io_cpu_s2_xcpt_pf_ld,
  output        io_cpu_s2_xcpt_pf_st,
  output        io_cpu_s2_xcpt_ae_ld,
  output        io_cpu_s2_xcpt_ae_st,
  output        io_cpu_ordered,
  output        io_cpu_perf_grant,
  input         io_cpu_keep_clock_enabled,
  output        io_cpu_clock_enabled,
  input         io_ptw_req_ready,
  output        io_ptw_req_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  input         io_ptw_resp_valid,
  input         io_ptw_resp_bits_ae,
  input  [53:0] io_ptw_resp_bits_pte_ppn,
  input         io_ptw_resp_bits_pte_d,
  input         io_ptw_resp_bits_pte_a,
  input         io_ptw_resp_bits_pte_g,
  input         io_ptw_resp_bits_pte_u,
  input         io_ptw_resp_bits_pte_x,
  input         io_ptw_resp_bits_pte_w,
  input         io_ptw_resp_bits_pte_r,
  input         io_ptw_resp_bits_pte_v,
  input  [1:0]  io_ptw_resp_bits_level,
  input         io_ptw_resp_bits_homogeneous,
  input  [3:0]  io_ptw_ptbr_mode,
  input  [1:0]  io_ptw_status_dprv,
  input         io_ptw_status_mxr,
  input         io_ptw_status_sum,
  input         io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
  input         io_ptw_pmp_0_cfg_w,
  input         io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr,
  input  [31:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
  input         io_ptw_pmp_1_cfg_w,
  input         io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr,
  input  [31:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
  input         io_ptw_pmp_2_cfg_w,
  input         io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr,
  input  [31:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
  input         io_ptw_pmp_3_cfg_w,
  input         io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr,
  input  [31:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
  input         io_ptw_pmp_4_cfg_w,
  input         io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr,
  input  [31:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
  input         io_ptw_pmp_5_cfg_w,
  input         io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr,
  input  [31:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
  input         io_ptw_pmp_6_cfg_w,
  input         io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr,
  input  [31:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
  input         io_ptw_pmp_7_cfg_w,
  input         io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr,
  input  [31:0] io_ptw_pmp_7_mask,
  input  [26:0] io_ptw_vpoffset_bits_value,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         data_halt,
  input         tlb_halt
);
  wire  metaArb_io_in_0_valid; // @[DCache.scala 98:23]
  wire [39:0] metaArb_io_in_0_bits_addr; // @[DCache.scala 98:23]
  wire [5:0] metaArb_io_in_0_bits_idx; // @[DCache.scala 98:23]
  wire [21:0] metaArb_io_in_0_bits_data; // @[DCache.scala 98:23]
  wire  metaArb_io_in_2_valid; // @[DCache.scala 98:23]
  wire [39:0] metaArb_io_in_2_bits_addr; // @[DCache.scala 98:23]
  wire [5:0] metaArb_io_in_2_bits_idx; // @[DCache.scala 98:23]
  wire [3:0] metaArb_io_in_2_bits_way_en; // @[DCache.scala 98:23]
  wire [21:0] metaArb_io_in_2_bits_data; // @[DCache.scala 98:23]
  wire  metaArb_io_in_3_valid; // @[DCache.scala 98:23]
  wire [39:0] metaArb_io_in_3_bits_addr; // @[DCache.scala 98:23]
  wire [5:0] metaArb_io_in_3_bits_idx; // @[DCache.scala 98:23]
  wire [3:0] metaArb_io_in_3_bits_way_en; // @[DCache.scala 98:23]
  wire [21:0] metaArb_io_in_3_bits_data; // @[DCache.scala 98:23]
  wire  metaArb_io_in_4_ready; // @[DCache.scala 98:23]
  wire  metaArb_io_in_4_valid; // @[DCache.scala 98:23]
  wire [39:0] metaArb_io_in_4_bits_addr; // @[DCache.scala 98:23]
  wire [5:0] metaArb_io_in_4_bits_idx; // @[DCache.scala 98:23]
  wire [3:0] metaArb_io_in_4_bits_way_en; // @[DCache.scala 98:23]
  wire [21:0] metaArb_io_in_4_bits_data; // @[DCache.scala 98:23]
  wire  metaArb_io_in_5_ready; // @[DCache.scala 98:23]
  wire  metaArb_io_in_5_valid; // @[DCache.scala 98:23]
  wire [39:0] metaArb_io_in_5_bits_addr; // @[DCache.scala 98:23]
  wire [5:0] metaArb_io_in_5_bits_idx; // @[DCache.scala 98:23]
  wire [3:0] metaArb_io_in_5_bits_way_en; // @[DCache.scala 98:23]
  wire [21:0] metaArb_io_in_5_bits_data; // @[DCache.scala 98:23]
  wire  metaArb_io_in_6_ready; // @[DCache.scala 98:23]
  wire  metaArb_io_in_6_valid; // @[DCache.scala 98:23]
  wire [39:0] metaArb_io_in_6_bits_addr; // @[DCache.scala 98:23]
  wire [5:0] metaArb_io_in_6_bits_idx; // @[DCache.scala 98:23]
  wire [3:0] metaArb_io_in_6_bits_way_en; // @[DCache.scala 98:23]
  wire [21:0] metaArb_io_in_6_bits_data; // @[DCache.scala 98:23]
  wire  metaArb_io_in_7_ready; // @[DCache.scala 98:23]
  wire  metaArb_io_in_7_valid; // @[DCache.scala 98:23]
  wire [39:0] metaArb_io_in_7_bits_addr; // @[DCache.scala 98:23]
  wire [5:0] metaArb_io_in_7_bits_idx; // @[DCache.scala 98:23]
  wire [3:0] metaArb_io_in_7_bits_way_en; // @[DCache.scala 98:23]
  wire [21:0] metaArb_io_in_7_bits_data; // @[DCache.scala 98:23]
  wire  metaArb_io_out_ready; // @[DCache.scala 98:23]
  wire  metaArb_io_out_valid; // @[DCache.scala 98:23]
  wire  metaArb_io_out_bits_write; // @[DCache.scala 98:23]
  wire [39:0] metaArb_io_out_bits_addr; // @[DCache.scala 98:23]
  wire [5:0] metaArb_io_out_bits_idx; // @[DCache.scala 98:23]
  wire [3:0] metaArb_io_out_bits_way_en; // @[DCache.scala 98:23]
  wire [21:0] metaArb_io_out_bits_data; // @[DCache.scala 98:23]
  wire [29:0] metaArb_io_covSum; // @[DCache.scala 98:23]
  wire  metaArb_metaAssert; // @[DCache.scala 98:23]
  reg [21:0] tag_array_0 [0:63]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_0;
  wire [21:0] tag_array_0_s1_meta_data; // @[DescribedSRAM.scala 23:21]
  wire [5:0] tag_array_0_s1_meta_addr; // @[DescribedSRAM.scala 23:21]
  wire [21:0] tag_array_0__T_567_data; // @[DescribedSRAM.scala 23:21]
  wire [5:0] tag_array_0__T_567_addr; // @[DescribedSRAM.scala 23:21]
  wire  tag_array_0__T_567_mask; // @[DescribedSRAM.scala 23:21]
  wire  tag_array_0__T_567_en; // @[DescribedSRAM.scala 23:21]
  reg  tag_array_0_s1_meta_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [5:0] tag_array_0_s1_meta_addr_pipe_0;
  reg [31:0] _RAND_2;
  reg [21:0] tag_array_1 [0:63]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_3;
  wire [21:0] tag_array_1_s1_meta_data; // @[DescribedSRAM.scala 23:21]
  wire [5:0] tag_array_1_s1_meta_addr; // @[DescribedSRAM.scala 23:21]
  wire [21:0] tag_array_1__T_567_data; // @[DescribedSRAM.scala 23:21]
  wire [5:0] tag_array_1__T_567_addr; // @[DescribedSRAM.scala 23:21]
  wire  tag_array_1__T_567_mask; // @[DescribedSRAM.scala 23:21]
  wire  tag_array_1__T_567_en; // @[DescribedSRAM.scala 23:21]
  reg  tag_array_1_s1_meta_en_pipe_0;
  reg [31:0] _RAND_4;
  reg [5:0] tag_array_1_s1_meta_addr_pipe_0;
  reg [31:0] _RAND_5;
  reg [21:0] tag_array_2 [0:63]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_6;
  wire [21:0] tag_array_2_s1_meta_data; // @[DescribedSRAM.scala 23:21]
  wire [5:0] tag_array_2_s1_meta_addr; // @[DescribedSRAM.scala 23:21]
  wire [21:0] tag_array_2__T_567_data; // @[DescribedSRAM.scala 23:21]
  wire [5:0] tag_array_2__T_567_addr; // @[DescribedSRAM.scala 23:21]
  wire  tag_array_2__T_567_mask; // @[DescribedSRAM.scala 23:21]
  wire  tag_array_2__T_567_en; // @[DescribedSRAM.scala 23:21]
  reg  tag_array_2_s1_meta_en_pipe_0;
  reg [31:0] _RAND_7;
  reg [5:0] tag_array_2_s1_meta_addr_pipe_0;
  reg [31:0] _RAND_8;
  reg [21:0] tag_array_3 [0:63]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_9;
  wire [21:0] tag_array_3_s1_meta_data; // @[DescribedSRAM.scala 23:21]
  wire [5:0] tag_array_3_s1_meta_addr; // @[DescribedSRAM.scala 23:21]
  wire [21:0] tag_array_3__T_567_data; // @[DescribedSRAM.scala 23:21]
  wire [5:0] tag_array_3__T_567_addr; // @[DescribedSRAM.scala 23:21]
  wire  tag_array_3__T_567_mask; // @[DescribedSRAM.scala 23:21]
  wire  tag_array_3__T_567_en; // @[DescribedSRAM.scala 23:21]
  reg  tag_array_3_s1_meta_en_pipe_0;
  reg [31:0] _RAND_10;
  reg [5:0] tag_array_3_s1_meta_addr_pipe_0;
  reg [31:0] _RAND_11;
  wire  data_clock; // @[DCache.scala 108:20]
  wire  data_io_req_valid; // @[DCache.scala 108:20]
  wire [11:0] data_io_req_bits_addr; // @[DCache.scala 108:20]
  wire  data_io_req_bits_write; // @[DCache.scala 108:20]
  wire [63:0] data_io_req_bits_wdata; // @[DCache.scala 108:20]
  wire [7:0] data_io_req_bits_eccMask; // @[DCache.scala 108:20]
  wire [3:0] data_io_req_bits_way_en; // @[DCache.scala 108:20]
  wire [63:0] data_io_resp_0; // @[DCache.scala 108:20]
  wire [63:0] data_io_resp_1; // @[DCache.scala 108:20]
  wire [63:0] data_io_resp_2; // @[DCache.scala 108:20]
  wire [63:0] data_io_resp_3; // @[DCache.scala 108:20]
  wire [29:0] data_io_covSum; // @[DCache.scala 108:20]
  wire  data_metaAssert; // @[DCache.scala 108:20]
  wire  data_metaReset; // @[DCache.scala 108:20]
  wire  dataArb_io_in_0_valid; // @[DCache.scala 109:23]
  wire [11:0] dataArb_io_in_0_bits_addr; // @[DCache.scala 109:23]
  wire  dataArb_io_in_0_bits_write; // @[DCache.scala 109:23]
  wire [63:0] dataArb_io_in_0_bits_wdata; // @[DCache.scala 109:23]
  wire [7:0] dataArb_io_in_0_bits_eccMask; // @[DCache.scala 109:23]
  wire [3:0] dataArb_io_in_0_bits_way_en; // @[DCache.scala 109:23]
  wire  dataArb_io_in_1_ready; // @[DCache.scala 109:23]
  wire  dataArb_io_in_1_valid; // @[DCache.scala 109:23]
  wire [11:0] dataArb_io_in_1_bits_addr; // @[DCache.scala 109:23]
  wire  dataArb_io_in_1_bits_write; // @[DCache.scala 109:23]
  wire [63:0] dataArb_io_in_1_bits_wdata; // @[DCache.scala 109:23]
  wire [7:0] dataArb_io_in_1_bits_eccMask; // @[DCache.scala 109:23]
  wire [3:0] dataArb_io_in_1_bits_way_en; // @[DCache.scala 109:23]
  wire  dataArb_io_in_2_ready; // @[DCache.scala 109:23]
  wire  dataArb_io_in_2_valid; // @[DCache.scala 109:23]
  wire [11:0] dataArb_io_in_2_bits_addr; // @[DCache.scala 109:23]
  wire [63:0] dataArb_io_in_2_bits_wdata; // @[DCache.scala 109:23]
  wire [7:0] dataArb_io_in_2_bits_eccMask; // @[DCache.scala 109:23]
  wire  dataArb_io_in_3_ready; // @[DCache.scala 109:23]
  wire  dataArb_io_in_3_valid; // @[DCache.scala 109:23]
  wire [11:0] dataArb_io_in_3_bits_addr; // @[DCache.scala 109:23]
  wire [63:0] dataArb_io_in_3_bits_wdata; // @[DCache.scala 109:23]
  wire [7:0] dataArb_io_in_3_bits_eccMask; // @[DCache.scala 109:23]
  wire  dataArb_io_out_valid; // @[DCache.scala 109:23]
  wire [11:0] dataArb_io_out_bits_addr; // @[DCache.scala 109:23]
  wire  dataArb_io_out_bits_write; // @[DCache.scala 109:23]
  wire [63:0] dataArb_io_out_bits_wdata; // @[DCache.scala 109:23]
  wire [7:0] dataArb_io_out_bits_eccMask; // @[DCache.scala 109:23]
  wire [3:0] dataArb_io_out_bits_way_en; // @[DCache.scala 109:23]
  wire [29:0] dataArb_io_covSum; // @[DCache.scala 109:23]
  wire  dataArb_metaAssert; // @[DCache.scala 109:23]
  wire  tlb_clock; // @[DCache.scala 184:19]
  wire  tlb_reset; // @[DCache.scala 184:19]
  wire  tlb_io_req_ready; // @[DCache.scala 184:19]
  wire  tlb_io_req_valid; // @[DCache.scala 184:19]
  wire [39:0] tlb_io_req_bits_vaddr; // @[DCache.scala 184:19]
  wire  tlb_io_req_bits_passthrough; // @[DCache.scala 184:19]
  wire [1:0] tlb_io_req_bits_size; // @[DCache.scala 184:19]
  wire [4:0] tlb_io_req_bits_cmd; // @[DCache.scala 184:19]
  wire  tlb_io_resp_miss; // @[DCache.scala 184:19]
  wire [31:0] tlb_io_resp_paddr; // @[DCache.scala 184:19]
  wire  tlb_io_resp_pf_ld; // @[DCache.scala 184:19]
  wire  tlb_io_resp_pf_st; // @[DCache.scala 184:19]
  wire  tlb_io_resp_ae_ld; // @[DCache.scala 184:19]
  wire  tlb_io_resp_ae_st; // @[DCache.scala 184:19]
  wire  tlb_io_resp_ma_ld; // @[DCache.scala 184:19]
  wire  tlb_io_resp_ma_st; // @[DCache.scala 184:19]
  wire  tlb_io_resp_cacheable; // @[DCache.scala 184:19]
  wire  tlb_io_sfence_valid; // @[DCache.scala 184:19]
  wire  tlb_io_sfence_bits_rs1; // @[DCache.scala 184:19]
  wire  tlb_io_sfence_bits_rs2; // @[DCache.scala 184:19]
  wire [38:0] tlb_io_sfence_bits_addr; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_req_ready; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_req_valid; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_req_bits_valid; // @[DCache.scala 184:19]
  wire [26:0] tlb_io_ptw_req_bits_bits_addr; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_resp_valid; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_resp_bits_ae; // @[DCache.scala 184:19]
  wire [53:0] tlb_io_ptw_resp_bits_pte_ppn; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_resp_bits_pte_d; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_resp_bits_pte_a; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_resp_bits_pte_g; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_resp_bits_pte_u; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_resp_bits_pte_x; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_resp_bits_pte_w; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_resp_bits_pte_r; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_resp_bits_pte_v; // @[DCache.scala 184:19]
  wire [1:0] tlb_io_ptw_resp_bits_level; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_resp_bits_homogeneous; // @[DCache.scala 184:19]
  wire [3:0] tlb_io_ptw_ptbr_mode; // @[DCache.scala 184:19]
  wire [1:0] tlb_io_ptw_status_dprv; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_status_mxr; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_status_sum; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_0_cfg_l; // @[DCache.scala 184:19]
  wire [1:0] tlb_io_ptw_pmp_0_cfg_a; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_0_cfg_x; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_0_cfg_w; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_0_cfg_r; // @[DCache.scala 184:19]
  wire [29:0] tlb_io_ptw_pmp_0_addr; // @[DCache.scala 184:19]
  wire [31:0] tlb_io_ptw_pmp_0_mask; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_1_cfg_l; // @[DCache.scala 184:19]
  wire [1:0] tlb_io_ptw_pmp_1_cfg_a; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_1_cfg_x; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_1_cfg_w; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_1_cfg_r; // @[DCache.scala 184:19]
  wire [29:0] tlb_io_ptw_pmp_1_addr; // @[DCache.scala 184:19]
  wire [31:0] tlb_io_ptw_pmp_1_mask; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_2_cfg_l; // @[DCache.scala 184:19]
  wire [1:0] tlb_io_ptw_pmp_2_cfg_a; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_2_cfg_x; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_2_cfg_w; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_2_cfg_r; // @[DCache.scala 184:19]
  wire [29:0] tlb_io_ptw_pmp_2_addr; // @[DCache.scala 184:19]
  wire [31:0] tlb_io_ptw_pmp_2_mask; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_3_cfg_l; // @[DCache.scala 184:19]
  wire [1:0] tlb_io_ptw_pmp_3_cfg_a; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_3_cfg_x; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_3_cfg_w; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_3_cfg_r; // @[DCache.scala 184:19]
  wire [29:0] tlb_io_ptw_pmp_3_addr; // @[DCache.scala 184:19]
  wire [31:0] tlb_io_ptw_pmp_3_mask; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_4_cfg_l; // @[DCache.scala 184:19]
  wire [1:0] tlb_io_ptw_pmp_4_cfg_a; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_4_cfg_x; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_4_cfg_w; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_4_cfg_r; // @[DCache.scala 184:19]
  wire [29:0] tlb_io_ptw_pmp_4_addr; // @[DCache.scala 184:19]
  wire [31:0] tlb_io_ptw_pmp_4_mask; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_5_cfg_l; // @[DCache.scala 184:19]
  wire [1:0] tlb_io_ptw_pmp_5_cfg_a; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_5_cfg_x; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_5_cfg_w; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_5_cfg_r; // @[DCache.scala 184:19]
  wire [29:0] tlb_io_ptw_pmp_5_addr; // @[DCache.scala 184:19]
  wire [31:0] tlb_io_ptw_pmp_5_mask; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_6_cfg_l; // @[DCache.scala 184:19]
  wire [1:0] tlb_io_ptw_pmp_6_cfg_a; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_6_cfg_x; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_6_cfg_w; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_6_cfg_r; // @[DCache.scala 184:19]
  wire [29:0] tlb_io_ptw_pmp_6_addr; // @[DCache.scala 184:19]
  wire [31:0] tlb_io_ptw_pmp_6_mask; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_7_cfg_l; // @[DCache.scala 184:19]
  wire [1:0] tlb_io_ptw_pmp_7_cfg_a; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_7_cfg_x; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_7_cfg_w; // @[DCache.scala 184:19]
  wire  tlb_io_ptw_pmp_7_cfg_r; // @[DCache.scala 184:19]
  wire [29:0] tlb_io_ptw_pmp_7_addr; // @[DCache.scala 184:19]
  wire [31:0] tlb_io_ptw_pmp_7_mask; // @[DCache.scala 184:19]
  wire [26:0] tlb_io_ptw_vpoffset_bits_value; // @[DCache.scala 184:19]
  wire [29:0] tlb_io_covSum; // @[DCache.scala 184:19]
  wire  tlb_metaAssert; // @[DCache.scala 184:19]
  wire  tlb_metaReset; // @[DCache.scala 184:19]
  wire [7:0] amoalu_io_mask; // @[DCache.scala 743:24]
  wire [4:0] amoalu_io_cmd; // @[DCache.scala 743:24]
  wire [63:0] amoalu_io_lhs; // @[DCache.scala 743:24]
  wire [63:0] amoalu_io_rhs; // @[DCache.scala 743:24]
  wire [63:0] amoalu_io_out; // @[DCache.scala 743:24]
  wire [29:0] amoalu_io_covSum; // @[DCache.scala 743:24]
  wire  amoalu_metaAssert; // @[DCache.scala 743:24]
  reg  clock_en_reg; // @[DCache.scala 88:25]
  reg [31:0] _RAND_12;
  reg [15:0] lfsr; // @[LFSR.scala 22:23]
  reg [31:0] _RAND_13;
  wire  _T_251; // @[LFSR.scala 23:43]
  wire  _T_253; // @[LFSR.scala 23:51]
  wire  _T_255; // @[LFSR.scala 23:59]
  wire [15:0] _T_257; // @[Cat.scala 30:58]
  wire  grantIsUncachedData; // @[package.scala 14:47]
  reg  blockUncachedGrant; // @[DCache.scala 572:31]
  reg [31:0] _RAND_14;
  reg  s1_valid; // @[DCache.scala 131:21]
  reg [31:0] _RAND_15;
  wire  _T_3218; // @[DCache.scala 574:52]
  wire  _T_3219; // @[DCache.scala 574:29]
  wire  grantIsRefill; // @[DCache.scala 491:29]
  wire  _T_3130; // @[DCache.scala 544:23]
  wire  _T_3082; // @[package.scala 14:47]
  wire  grantIsCached; // @[package.scala 14:62]
  reg [8:0] _T_3069; // @[Edges.scala 229:27]
  reg [31:0] _RAND_16;
  wire  d_first; // @[Edges.scala 231:25]
  wire  _T_3091; // @[DCache.scala 496:50]
  wire  _T_3093; // @[DCache.scala 496:24]
  wire  _GEN_169; // @[DCache.scala 544:51]
  wire  tl_out__d_ready; // @[DCache.scala 574:66]
  wire  _T_3094; // @[Decoupled.scala 37:37]
  wire  _T_3073; // @[Edges.scala 232:25]
  wire [26:0] _T_3062; // @[package.scala 185:77]
  wire [8:0] _T_3065; // @[Edges.scala 220:59]
  wire [8:0] _T_3067; // @[Edges.scala 221:14]
  wire  _T_3074; // @[Edges.scala 232:47]
  wire  d_last; // @[Edges.scala 232:37]
  wire  _GEN_147; // @[DCache.scala 498:26]
  wire  _GEN_159; // @[DCache.scala 497:26]
  wire [63:0] _T_270; // @[DCache.scala 112:65]
  wire [31:0] _T_281; // @[Cat.scala 30:58]
  wire [31:0] _T_284; // @[Cat.scala 30:58]
  wire  _T_288; // @[Decoupled.scala 37:37]
  reg  s1_probe; // @[DCache.scala 132:21]
  reg [31:0] _RAND_17;
  reg  s2_probe; // @[DCache.scala 232:21]
  reg [31:0] _RAND_18;
  wire  _T_734; // @[DCache.scala 233:34]
  reg [2:0] release_state; // @[DCache.scala 155:26]
  reg [31:0] _RAND_19;
  wire  _T_735; // @[DCache.scala 233:63]
  wire  releaseInFlight; // @[DCache.scala 233:46]
  reg  grantInProgress; // @[DCache.scala 492:28]
  reg [31:0] _RAND_20;
  wire  _T_3223; // @[DCache.scala 587:37]
  reg [2:0] blockProbeAfterGrantCount; // @[DCache.scala 493:38]
  reg [31:0] _RAND_21;
  wire  _T_3224; // @[DCache.scala 587:85]
  wire  _T_3225; // @[DCache.scala 587:56]
  reg [6:0] lrscCount; // @[DCache.scala 327:22]
  reg [31:0] _RAND_22;
  wire  lrscValid; // @[DCache.scala 328:29]
  wire  block_probe; // @[DCache.scala 587:89]
  wire  _T_3230; // @[DCache.scala 589:44]
  wire  _T_3232; // @[DCache.scala 589:60]
  reg  s2_valid_pre_xcpt; // @[DCache.scala 230:30]
  reg [31:0] _RAND_23;
  wire [5:0] _T_730; // @[DCache.scala 231:55]
  wire  _T_731; // @[DCache.scala 231:62]
  wire  s2_valid; // @[DCache.scala 231:36]
  wire  tl_out__b_ready; // @[DCache.scala 589:73]
  wire  _T_290; // @[Decoupled.scala 37:37]
  reg [1:0] probe_bits_param; // @[Reg.scala 11:16]
  reg [31:0] _RAND_24;
  reg [3:0] probe_bits_size; // @[Reg.scala 11:16]
  reg [31:0] _RAND_25;
  reg  probe_bits_source; // @[Reg.scala 11:16]
  reg [31:0] _RAND_26;
  reg [31:0] probe_bits_address; // @[Reg.scala 11:16]
  reg [31:0] _RAND_27;
  wire  s1_valid_masked; // @[DCache.scala 135:34]
  reg [1:0] s2_probe_state_state; // @[Reg.scala 11:16]
  reg [31:0] _RAND_28;
  wire [3:0] _T_1069; // @[Cat.scala 30:58]
  wire  _T_1126; // @[Misc.scala 58:20]
  wire  _T_1122; // @[Misc.scala 58:20]
  wire  _T_1118; // @[Misc.scala 58:20]
  wire  _T_1114; // @[Misc.scala 58:20]
  wire  _T_1110; // @[Misc.scala 58:20]
  wire  _T_1106; // @[Misc.scala 58:20]
  wire  _T_1102; // @[Misc.scala 58:20]
  wire  _T_1098; // @[Misc.scala 58:20]
  wire  _T_1094; // @[Misc.scala 58:20]
  wire  _T_1090; // @[Misc.scala 58:20]
  wire  _T_1086; // @[Misc.scala 58:20]
  wire  _T_1082; // @[Misc.scala 58:20]
  wire  _T_1099; // @[Misc.scala 40:9]
  wire  _T_1103; // @[Misc.scala 40:9]
  wire  _T_1107; // @[Misc.scala 40:9]
  wire  _T_1111; // @[Misc.scala 40:9]
  wire  _T_1115; // @[Misc.scala 40:9]
  wire  _T_1119; // @[Misc.scala 40:9]
  wire  _T_1123; // @[Misc.scala 40:9]
  wire  s2_prb_ack_data; // @[Misc.scala 40:9]
  wire  _T_3304; // @[Metadata.scala 50:45]
  reg [8:0] _T_3247; // @[Edges.scala 229:27]
  reg [31:0] _RAND_29;
  wire  _T_3251; // @[Edges.scala 232:25]
  wire  _T_3315; // @[package.scala 14:47]
  wire  _T_3316; // @[package.scala 14:47]
  wire  _T_3317; // @[package.scala 14:62]
  wire  _T_3314; // @[DCache.scala 655:25]
  wire  _T_3313; // @[DCache.scala 650:25]
  wire [2:0] _GEN_251; // @[DCache.scala 655:48]
  wire [2:0] tl_out__c_bits_opcode; // @[DCache.scala 659:81]
  wire [3:0] tl_out__c_bits_size; // @[DCache.scala 659:81]
  wire [26:0] _T_3240; // @[package.scala 185:77]
  wire [8:0] _T_3243; // @[Edges.scala 220:59]
  wire [8:0] _T_3245; // @[Edges.scala 221:14]
  wire  _T_3252; // @[Edges.scala 232:47]
  wire  c_last; // @[Edges.scala 232:37]
  wire  _T_3312; // @[DCache.scala 646:25]
  reg  s2_release_data_valid; // @[DCache.scala 600:34]
  reg [31:0] _RAND_30;
  wire  _GEN_200; // @[DCache.scala 624:36]
  wire  _GEN_221; // @[DCache.scala 620:21]
  wire  _GEN_238; // @[DCache.scala 646:47]
  wire  tl_out__c_valid; // @[DCache.scala 650:48]
  wire  _T_3238; // @[Decoupled.scala 37:37]
  wire  releaseDone; // @[Edges.scala 233:22]
  wire  _GEN_198; // @[DCache.scala 626:45]
  wire  probeNack; // @[DCache.scala 624:36]
  reg [4:0] s1_req_cmd; // @[DCache.scala 137:19]
  reg [31:0] _RAND_31;
  wire  _T_302; // @[Consts.scala 93:31]
  wire  _T_303; // @[Consts.scala 93:48]
  wire  _T_304; // @[Consts.scala 93:41]
  wire  _T_305; // @[Consts.scala 93:65]
  wire  _T_306; // @[Consts.scala 93:58]
  wire  _T_307; // @[package.scala 14:47]
  wire  _T_308; // @[package.scala 14:47]
  wire  _T_311; // @[package.scala 14:62]
  wire  _T_309; // @[package.scala 14:47]
  wire  _T_312; // @[package.scala 14:62]
  wire  _T_310; // @[package.scala 14:47]
  wire  _T_313; // @[package.scala 14:62]
  wire  _T_314; // @[package.scala 14:47]
  wire  _T_315; // @[package.scala 14:47]
  wire  _T_319; // @[package.scala 14:62]
  wire  _T_316; // @[package.scala 14:47]
  wire  _T_320; // @[package.scala 14:62]
  wire  _T_317; // @[package.scala 14:47]
  wire  _T_321; // @[package.scala 14:62]
  wire  _T_318; // @[package.scala 14:47]
  wire  _T_322; // @[package.scala 14:62]
  wire  _T_323; // @[Consts.scala 91:44]
  wire  s1_read; // @[Consts.scala 93:75]
  reg  _T_738; // @[DCache.scala 234:40]
  reg [31:0] _RAND_32;
  wire  s2_valid_masked; // @[DCache.scala 234:34]
  reg [4:0] s2_req_cmd; // @[DCache.scala 236:19]
  reg [31:0] _RAND_33;
  wire  _T_749; // @[Consts.scala 93:31]
  wire  _T_750; // @[Consts.scala 93:48]
  wire  _T_751; // @[Consts.scala 93:41]
  wire  _T_752; // @[Consts.scala 93:65]
  wire  _T_753; // @[Consts.scala 93:58]
  wire  _T_754; // @[package.scala 14:47]
  wire  _T_755; // @[package.scala 14:47]
  wire  _T_758; // @[package.scala 14:62]
  wire  _T_756; // @[package.scala 14:47]
  wire  _T_759; // @[package.scala 14:62]
  wire  _T_757; // @[package.scala 14:47]
  wire  _T_760; // @[package.scala 14:62]
  wire  _T_761; // @[package.scala 14:47]
  wire  _T_762; // @[package.scala 14:47]
  wire  _T_766; // @[package.scala 14:62]
  wire  _T_763; // @[package.scala 14:47]
  wire  _T_767; // @[package.scala 14:62]
  wire  _T_764; // @[package.scala 14:47]
  wire  _T_768; // @[package.scala 14:62]
  wire  _T_765; // @[package.scala 14:47]
  wire  _T_769; // @[package.scala 14:62]
  wire  _T_770; // @[Consts.scala 91:44]
  wire  s2_read; // @[Consts.scala 93:75]
  wire  _T_771; // @[Consts.scala 94:32]
  wire  _T_772; // @[Consts.scala 94:49]
  wire  _T_773; // @[Consts.scala 94:42]
  wire  _T_775; // @[Consts.scala 94:59]
  wire  s2_write; // @[Consts.scala 94:76]
  wire  s2_readwrite; // @[DCache.scala 247:30]
  wire  _T_1033; // @[DCache.scala 282:51]
  wire  _T_926; // @[Consts.scala 95:54]
  wire  _T_927; // @[Consts.scala 95:47]
  wire  _T_929; // @[Consts.scala 95:64]
  reg [1:0] s2_hit_state_state; // @[Reg.scala 11:16]
  reg [31:0] _RAND_34;
  wire [3:0] _T_931; // @[Cat.scala 30:58]
  wire  _T_989; // @[Misc.scala 51:20]
  wire  _T_986; // @[Misc.scala 51:20]
  wire  _T_983; // @[Misc.scala 51:20]
  wire  _T_980; // @[Misc.scala 51:20]
  wire  _T_977; // @[Misc.scala 51:20]
  wire  _T_974; // @[Misc.scala 51:20]
  wire  _T_971; // @[Misc.scala 51:20]
  wire  _T_968; // @[Misc.scala 51:20]
  wire  _T_965; // @[Misc.scala 51:20]
  wire  _T_962; // @[Misc.scala 51:20]
  wire  _T_959; // @[Misc.scala 51:20]
  wire  _T_956; // @[Misc.scala 51:20]
  wire  _T_975; // @[Misc.scala 37:9]
  wire  _T_978; // @[Misc.scala 37:9]
  wire  _T_981; // @[Misc.scala 37:9]
  wire  _T_984; // @[Misc.scala 37:9]
  wire  _T_987; // @[Misc.scala 37:9]
  wire  s2_hit; // @[Misc.scala 37:9]
  wire  s2_valid_hit_pre_data_ecc; // @[DCache.scala 282:85]
  wire  _T_1417; // @[DCache.scala 345:46]
  reg [33:0] lrscAddr; // @[DCache.scala 330:21]
  reg [63:0] _RAND_35;
  reg [39:0] s2_req_addr; // @[DCache.scala 236:19]
  reg [63:0] _RAND_36;
  wire  lrscAddrMatch; // @[DCache.scala 331:32]
  wire  _T_1255; // @[DCache.scala 332:41]
  wire  s2_sc_fail; // @[DCache.scala 332:26]
  wire  _T_1419; // @[DCache.scala 345:58]
  reg  pstore1_held; // @[DCache.scala 359:25]
  reg [31:0] _RAND_37;
  wire  pstore1_valid_pre_kill; // @[DCache.scala 361:56]
  reg [39:0] pstore1_addr; // @[Reg.scala 11:16]
  reg [63:0] _RAND_38;
  reg [39:0] s1_req_addr; // @[DCache.scala 137:19]
  reg [63:0] _RAND_39;
  wire  _T_1591; // @[DCache.scala 414:31]
  wire  _T_324; // @[Consts.scala 94:32]
  wire  _T_325; // @[Consts.scala 94:49]
  wire  _T_326; // @[Consts.scala 94:42]
  wire  _T_328; // @[Consts.scala 94:59]
  wire  s1_write; // @[Consts.scala 94:76]
  reg [7:0] pstore1_mask; // @[Reg.scala 11:16]
  reg [31:0] _RAND_40;
  wire [7:0] _T_1614; // @[Cat.scala 30:58]
  wire [7:0] _T_1629; // @[Cat.scala 30:58]
  reg [2:0] s1_req_typ; // @[DCache.scala 137:19]
  reg [31:0] _RAND_41;
  wire  _T_701; // @[AMOALU.scala 17:57]
  wire  _T_703; // @[AMOALU.scala 17:46]
  wire  _T_705; // @[AMOALU.scala 18:22]
  wire [1:0] _T_706; // @[Cat.scala 30:58]
  wire [1:0] _T_708; // @[AMOALU.scala 17:22]
  wire  _T_709; // @[AMOALU.scala 17:57]
  wire [1:0] _T_710; // @[AMOALU.scala 17:51]
  wire [1:0] _T_711; // @[AMOALU.scala 17:46]
  wire [1:0] _T_713; // @[AMOALU.scala 18:22]
  wire [3:0] _T_714; // @[Cat.scala 30:58]
  wire [3:0] _T_716; // @[AMOALU.scala 17:22]
  wire  _T_717; // @[AMOALU.scala 17:57]
  wire [3:0] _T_718; // @[AMOALU.scala 17:51]
  wire [3:0] _T_719; // @[AMOALU.scala 17:46]
  wire [3:0] _T_721; // @[AMOALU.scala 18:22]
  wire [7:0] _T_722; // @[Cat.scala 30:58]
  wire [7:0] s1_mask; // @[DCache.scala 228:20]
  wire [7:0] _T_1652; // @[Cat.scala 30:58]
  wire [7:0] _T_1667; // @[Cat.scala 30:58]
  wire [7:0] _T_1668; // @[DCache.scala 415:38]
  wire  _T_1669; // @[DCache.scala 415:62]
  wire [7:0] _T_1670; // @[DCache.scala 415:73]
  wire  _T_1671; // @[DCache.scala 415:84]
  wire  _T_1672; // @[DCache.scala 415:8]
  wire  _T_1673; // @[DCache.scala 414:68]
  wire  _T_1674; // @[DCache.scala 417:29]
  reg  pstore2_valid; // @[DCache.scala 356:26]
  reg [31:0] _RAND_42;
  reg [39:0] pstore2_addr; // @[Reg.scala 11:16]
  reg [63:0] _RAND_43;
  wire  _T_1677; // @[DCache.scala 414:31]
  reg [7:0] mask; // @[DCache.scala 387:19]
  reg [31:0] _RAND_44;
  wire [7:0] _T_1700; // @[Cat.scala 30:58]
  wire [7:0] _T_1715; // @[Cat.scala 30:58]
  wire [7:0] _T_1754; // @[DCache.scala 415:38]
  wire  _T_1755; // @[DCache.scala 415:62]
  wire [7:0] _T_1756; // @[DCache.scala 415:73]
  wire  _T_1757; // @[DCache.scala 415:84]
  wire  _T_1758; // @[DCache.scala 415:8]
  wire  _T_1759; // @[DCache.scala 414:68]
  wire  _T_1760; // @[DCache.scala 418:21]
  wire  s1_hazard; // @[DCache.scala 417:71]
  wire  s1_raw_hazard; // @[DCache.scala 419:31]
  wire  _T_1761; // @[DCache.scala 424:18]
  wire [1:0] _T_958; // @[Misc.scala 37:36]
  wire [1:0] _T_961; // @[Misc.scala 37:36]
  wire [1:0] _T_964; // @[Misc.scala 37:36]
  wire [1:0] _T_967; // @[Misc.scala 37:36]
  wire [1:0] _T_970; // @[Misc.scala 37:36]
  wire [1:0] _T_973; // @[Misc.scala 37:36]
  wire [1:0] _T_976; // @[Misc.scala 37:36]
  wire [1:0] _T_979; // @[Misc.scala 37:36]
  wire [1:0] _T_982; // @[Misc.scala 37:36]
  wire [1:0] _T_985; // @[Misc.scala 37:36]
  wire [1:0] _T_988; // @[Misc.scala 37:36]
  wire [1:0] s2_grow_param; // @[Misc.scala 37:36]
  wire  _T_1195; // @[Metadata.scala 46:46]
  wire  s2_update_meta; // @[Metadata.scala 47:40]
  wire  _T_1201; // @[DCache.scala 301:41]
  wire  _T_1202; // @[DCache.scala 301:24]
  wire  s1_readwrite; // @[DCache.scala 146:30]
  wire  _T_543; // @[DCache.scala 193:18]
  wire  _T_544; // @[DCache.scala 193:34]
  wire  _GEN_74; // @[DCache.scala 301:61]
  wire  _GEN_98; // @[DCache.scala 424:36]
  wire  _GEN_219; // @[DCache.scala 635:24]
  wire  s1_nack; // @[DCache.scala 620:21]
  wire  s1_valid_not_nacked; // @[DCache.scala 136:38]
  reg [6:0] s1_req_tag; // @[DCache.scala 137:19]
  reg [31:0] _RAND_45;
  reg  s1_req_phys; // @[DCache.scala 137:19]
  reg [31:0] _RAND_46;
  wire  s0_clk_en; // @[DCache.scala 138:40]
  wire [39:0] _T_300; // @[Cat.scala 30:58]
  wire  _GEN_9; // @[DCache.scala 142:36]
  wire  s1_sfence; // @[DCache.scala 147:30]
  reg  s1_flush_valid; // @[DCache.scala 148:27]
  reg [31:0] _RAND_47;
  reg  cached_grant_wait; // @[DCache.scala 152:30]
  reg [31:0] _RAND_48;
  reg  release_ack_wait; // @[DCache.scala 153:29]
  reg [31:0] _RAND_49;
  wire  can_acquire_before_release; // @[DCache.scala 154:36]
  wire  inWriteback; // @[package.scala 14:62]
  wire  _T_357; // @[DCache.scala 159:38]
  wire  _T_359; // @[DCache.scala 159:51]
  wire  _T_361; // @[DCache.scala 159:73]
  reg  uncachedInFlight_0; // @[DCache.scala 162:33]
  reg [31:0] _RAND_50;
  reg [39:0] uncachedReqs_0_addr; // @[DCache.scala 163:25]
  reg [63:0] _RAND_51;
  reg [6:0] uncachedReqs_0_tag; // @[DCache.scala 163:25]
  reg [31:0] _RAND_52;
  reg [2:0] uncachedReqs_0_typ; // @[DCache.scala 163:25]
  reg [31:0] _RAND_53;
  wire  _T_388; // @[Consts.scala 93:31]
  wire  _T_389; // @[Consts.scala 93:48]
  wire  _T_390; // @[Consts.scala 93:41]
  wire  _T_391; // @[Consts.scala 93:65]
  wire  _T_392; // @[Consts.scala 93:58]
  wire  _T_393; // @[package.scala 14:47]
  wire  _T_394; // @[package.scala 14:47]
  wire  _T_395; // @[package.scala 14:47]
  wire  _T_396; // @[package.scala 14:47]
  wire  _T_397; // @[package.scala 14:62]
  wire  _T_398; // @[package.scala 14:62]
  wire  _T_399; // @[package.scala 14:62]
  wire  _T_400; // @[package.scala 14:47]
  wire  _T_401; // @[package.scala 14:47]
  wire  _T_402; // @[package.scala 14:47]
  wire  _T_403; // @[package.scala 14:47]
  wire  _T_404; // @[package.scala 14:47]
  wire  _T_405; // @[package.scala 14:62]
  wire  _T_406; // @[package.scala 14:62]
  wire  _T_407; // @[package.scala 14:62]
  wire  _T_408; // @[package.scala 14:62]
  wire  _T_409; // @[Consts.scala 91:44]
  wire  s0_read; // @[Consts.scala 93:75]
  wire  _T_410; // @[package.scala 14:47]
  wire  _T_411; // @[package.scala 14:47]
  wire  _T_412; // @[package.scala 14:62]
  wire  res; // @[DCache.scala 912:15]
  wire  _T_440; // @[Consts.scala 94:49]
  wire  _T_441; // @[Consts.scala 94:42]
  wire  _T_443; // @[Consts.scala 94:59]
  wire  _T_461; // @[Consts.scala 94:76]
  wire  _T_466; // @[DCache.scala 918:23]
  wire  _T_467; // @[DCache.scala 917:21]
  wire  _T_469; // @[DCache.scala 913:28]
  wire  _T_471; // @[DCache.scala 913:11]
  wire  _T_473; // @[DCache.scala 167:46]
  wire  _T_477; // @[DCache.scala 173:33]
  wire  _GEN_16; // @[DCache.scala 173:45]
  wire  _GEN_18; // @[DCache.scala 181:34]
  wire  _T_540; // @[DCache.scala 192:27]
  wire  _T_542; // @[DCache.scala 192:53]
  wire  _GEN_19; // @[DCache.scala 192:79]
  wire [1:0] s1_victim_way; // @[Replacement.scala 19:44]
  wire [21:0] _T_600;
  wire [21:0] _T_607;
  wire [21:0] _T_614;
  wire [21:0] _T_621;
  wire [19:0] s1_tag; // @[DCache.scala 219:29]
  wire  _T_624; // @[Metadata.scala 50:45]
  wire  _T_625; // @[DCache.scala 220:83]
  wire  _T_626; // @[DCache.scala 220:74]
  wire  _T_627; // @[Metadata.scala 50:45]
  wire  _T_628; // @[DCache.scala 220:83]
  wire  _T_629; // @[DCache.scala 220:74]
  wire  _T_630; // @[Metadata.scala 50:45]
  wire  _T_631; // @[DCache.scala 220:83]
  wire  _T_632; // @[DCache.scala 220:74]
  wire  _T_633; // @[Metadata.scala 50:45]
  wire  _T_634; // @[DCache.scala 220:83]
  wire  _T_635; // @[DCache.scala 220:74]
  wire [3:0] s1_meta_hit_way; // @[Cat.scala 30:58]
  wire  _T_642; // @[DCache.scala 222:59]
  wire [1:0] _T_643; // @[DCache.scala 222:41]
  wire  _T_646; // @[DCache.scala 222:59]
  wire [1:0] _T_647; // @[DCache.scala 222:41]
  wire  _T_650; // @[DCache.scala 222:59]
  wire [1:0] _T_651; // @[DCache.scala 222:41]
  wire  _T_654; // @[DCache.scala 222:59]
  wire [1:0] _T_655; // @[DCache.scala 222:41]
  wire [1:0] _T_656; // @[DCache.scala 223:19]
  wire [1:0] _T_657; // @[DCache.scala 223:19]
  wire [1:0] s1_meta_hit_state_state; // @[DCache.scala 223:19]
  wire  _T_665; // @[package.scala 31:81]
  wire  _T_667; // @[package.scala 31:81]
  wire  _T_669; // @[package.scala 31:81]
  wire  s2_hit_valid; // @[Metadata.scala 50:45]
  reg [3:0] s2_hit_way; // @[Reg.scala 11:16]
  reg [31:0] _RAND_54;
  reg [1:0] _T_1060; // @[Reg.scala 11:16]
  reg [31:0] _RAND_55;
  wire [3:0] _T_1061; // @[OneHot.scala 45:35]
  wire [3:0] s2_victim_way; // @[DCache.scala 292:26]
  reg [3:0] s2_probe_way; // @[Reg.scala 11:16]
  reg [31:0] _RAND_56;
  wire [3:0] releaseWay; // @[DCache.scala 659:81]
  wire [3:0] _T_670; // @[DCache.scala 226:61]
  wire [63:0] s1_all_data_ways_4; // @[Cat.scala 30:58]
  wire  _T_724; // @[DCache.scala 230:52]
  reg [6:0] s2_req_tag; // @[DCache.scala 236:19]
  reg [31:0] _RAND_57;
  reg [2:0] s2_req_typ; // @[DCache.scala 236:19]
  reg [31:0] _RAND_58;
  reg  s2_uncached; // @[DCache.scala 237:24]
  reg [31:0] _RAND_59;
  wire  _T_742; // @[DCache.scala 239:29]
  reg [39:0] _T_746; // @[Reg.scala 11:16]
  reg [63:0] _RAND_60;
  wire [39:0] s2_vaddr; // @[Cat.scala 30:58]
  reg  s2_flush_valid_pre_tag_ecc; // @[DCache.scala 248:43]
  reg [31:0] _RAND_61;
  wire  en; // @[DCache.scala 258:23]
  wire  _T_3079; // @[package.scala 14:47]
  wire  _T_3081; // @[package.scala 14:62]
  wire  _T_3080; // @[package.scala 14:47]
  wire  grantIsUncached; // @[package.scala 14:62]
  wire [4:0] _GEN_129; // @[DCache.scala 516:34]
  wire [4:0] _GEN_137; // @[DCache.scala 507:35]
  wire [4:0] _GEN_149; // @[DCache.scala 498:26]
  wire [4:0] s1_data_way; // @[DCache.scala 497:26]
  wire [63:0] s1_all_data_ways_0; // @[DCache.scala 227:29 DCache.scala 227:29]
  wire [63:0] _T_859; // @[Mux.scala 19:72]
  wire [63:0] s1_all_data_ways_1; // @[DCache.scala 227:29 DCache.scala 227:29]
  wire [63:0] _T_860; // @[Mux.scala 19:72]
  wire [63:0] s1_all_data_ways_2; // @[DCache.scala 227:29 DCache.scala 227:29]
  wire [63:0] _T_861; // @[Mux.scala 19:72]
  wire [63:0] s1_all_data_ways_3; // @[DCache.scala 227:29 DCache.scala 227:29]
  wire [63:0] _T_862; // @[Mux.scala 19:72]
  wire [63:0] _T_863; // @[Mux.scala 19:72]
  wire [63:0] _T_864; // @[Mux.scala 19:72]
  wire [63:0] _T_865; // @[Mux.scala 19:72]
  wire [63:0] _T_866; // @[Mux.scala 19:72]
  wire [63:0] _T_867; // @[Mux.scala 19:72]
  wire  _T_871; // @[DCache.scala 264:58]
  reg [63:0] s2_data; // @[Reg.scala 11:16]
  reg [63:0] _RAND_62;
  wire [31:0] _T_1023; // @[Cat.scala 30:58]
  wire [31:0] _T_1026; // @[Cat.scala 30:58]
  wire [63:0] s2_data_corrected; // @[Cat.scala 30:58]
  wire  _T_1045; // @[DCache.scala 285:73]
  wire  s2_valid_miss; // @[DCache.scala 285:84]
  wire  _T_1047; // @[DCache.scala 286:44]
  wire  s2_valid_cached_miss; // @[DCache.scala 286:60]
  wire  s2_want_victimize; // @[DCache.scala 288:102]
  wire  _T_1054; // @[DCache.scala 291:49]
  wire  s2_valid_uncached_pending; // @[DCache.scala 291:64]
  reg [19:0] s2_victim_tag; // @[Reg.scala 11:16]
  reg [31:0] _RAND_63;
  reg [1:0] _T_1068_state; // @[Reg.scala 11:16]
  reg [31:0] _RAND_64;
  wire [1:0] s2_victim_state_state; // @[DCache.scala 294:28]
  wire [2:0] _T_1084; // @[Misc.scala 40:36]
  wire [2:0] _T_1088; // @[Misc.scala 40:36]
  wire [2:0] _T_1092; // @[Misc.scala 40:36]
  wire [2:0] _T_1096; // @[Misc.scala 40:36]
  wire [2:0] _T_1100; // @[Misc.scala 40:36]
  wire [2:0] _T_1104; // @[Misc.scala 40:36]
  wire [1:0] _T_1105; // @[Misc.scala 40:63]
  wire [2:0] _T_1108; // @[Misc.scala 40:36]
  wire [1:0] _T_1109; // @[Misc.scala 40:63]
  wire [2:0] _T_1112; // @[Misc.scala 40:36]
  wire [1:0] _T_1113; // @[Misc.scala 40:63]
  wire [2:0] _T_1116; // @[Misc.scala 40:36]
  wire [1:0] _T_1117; // @[Misc.scala 40:63]
  wire [2:0] _T_1120; // @[Misc.scala 40:36]
  wire [1:0] _T_1121; // @[Misc.scala 40:63]
  wire [2:0] _T_1124; // @[Misc.scala 40:36]
  wire [1:0] _T_1125; // @[Misc.scala 40:63]
  wire [2:0] s2_report_param; // @[Misc.scala 40:36]
  wire [1:0] probeNewCoh_state; // @[Misc.scala 40:63]
  wire [3:0] _T_1135; // @[Cat.scala 30:58]
  wire  _T_1148; // @[Misc.scala 58:20]
  wire [2:0] _T_1150; // @[Misc.scala 40:36]
  wire  _T_1152; // @[Misc.scala 58:20]
  wire [2:0] _T_1154; // @[Misc.scala 40:36]
  wire  _T_1156; // @[Misc.scala 58:20]
  wire [2:0] _T_1158; // @[Misc.scala 40:36]
  wire  _T_1160; // @[Misc.scala 58:20]
  wire [2:0] _T_1162; // @[Misc.scala 40:36]
  wire  _T_1164; // @[Misc.scala 58:20]
  wire  _T_1165; // @[Misc.scala 40:9]
  wire [2:0] _T_1166; // @[Misc.scala 40:36]
  wire  _T_1168; // @[Misc.scala 58:20]
  wire  _T_1169; // @[Misc.scala 40:9]
  wire [2:0] _T_1170; // @[Misc.scala 40:36]
  wire [1:0] _T_1171; // @[Misc.scala 40:63]
  wire  _T_1172; // @[Misc.scala 58:20]
  wire  _T_1173; // @[Misc.scala 40:9]
  wire [2:0] _T_1174; // @[Misc.scala 40:36]
  wire [1:0] _T_1175; // @[Misc.scala 40:63]
  wire  _T_1176; // @[Misc.scala 58:20]
  wire  _T_1177; // @[Misc.scala 40:9]
  wire [2:0] _T_1178; // @[Misc.scala 40:36]
  wire [1:0] _T_1179; // @[Misc.scala 40:63]
  wire  _T_1180; // @[Misc.scala 58:20]
  wire  _T_1181; // @[Misc.scala 40:9]
  wire [2:0] _T_1182; // @[Misc.scala 40:36]
  wire [1:0] _T_1183; // @[Misc.scala 40:63]
  wire  _T_1184; // @[Misc.scala 58:20]
  wire  _T_1185; // @[Misc.scala 40:9]
  wire [2:0] _T_1186; // @[Misc.scala 40:36]
  wire [1:0] _T_1187; // @[Misc.scala 40:63]
  wire  _T_1188; // @[Misc.scala 58:20]
  wire  _T_1189; // @[Misc.scala 40:9]
  wire [2:0] _T_1190; // @[Misc.scala 40:36]
  wire [1:0] _T_1191; // @[Misc.scala 40:63]
  wire  _T_1192; // @[Misc.scala 58:20]
  wire  s2_victim_dirty; // @[Misc.scala 40:9]
  wire [2:0] s2_shrink_param; // @[Misc.scala 40:36]
  wire [1:0] voluntaryNewCoh_state; // @[Misc.scala 40:63]
  wire  _T_1197; // @[DCache.scala 300:30]
  wire  _T_1198; // @[DCache.scala 300:78]
  wire  _T_1200; // @[DCache.scala 300:47]
  wire  _T_1234; // @[DCache.scala 317:84]
  wire [1:0] _T_1244_state; // @[DCache.scala 322:82]
  wire  _T_1251; // @[DCache.scala 329:34]
  wire  lrscBackingOff; // @[DCache.scala 329:38]
  wire  _T_1257; // @[DCache.scala 333:23]
  wire  _T_1259; // @[DCache.scala 333:32]
  wire  _T_1260; // @[DCache.scala 333:54]
  wire [6:0] _T_1268; // @[DCache.scala 337:49]
  wire  _T_1269; // @[DCache.scala 338:29]
  wire  _T_1278; // @[DCache.scala 347:63]
  reg [4:0] pstore1_cmd; // @[Reg.scala 11:16]
  reg [31:0] _RAND_65;
  reg [63:0] pstore1_data; // @[Reg.scala 11:16]
  reg [63:0] _RAND_66;
  reg [3:0] pstore1_way; // @[Reg.scala 11:16]
  reg [31:0] _RAND_67;
  wire  _T_1339; // @[DCache.scala 918:23]
  wire  _T_1340; // @[DCache.scala 917:21]
  reg  pstore1_rmw; // @[Reg.scala 11:16]
  reg [31:0] _RAND_68;
  wire  _T_1344; // @[DCache.scala 354:39]
  wire  pstore_drain_opportunistic; // @[DCache.scala 357:36]
  wire  pstore1_valid_likely; // @[DCache.scala 360:51]
  wire  _T_1426; // @[DCache.scala 365:54]
  wire  _T_1427; // @[DCache.scala 365:85]
  wire  _T_1428; // @[DCache.scala 365:98]
  wire  pstore_drain_structural; // @[DCache.scala 365:71]
  wire  _T_1438; // @[DCache.scala 366:63]
  wire  _T_1439; // @[DCache.scala 366:22]
  wire  _T_1441; // @[DCache.scala 366:9]
  wire  _T_1457; // @[DCache.scala 374:41]
  wire  _T_1458; // @[DCache.scala 374:58]
  wire  _T_1459; // @[DCache.scala 374:107]
  wire  _T_1460; // @[DCache.scala 374:76]
  wire  pstore_drain; // @[DCache.scala 373:48]
  wire  _T_1470; // @[DCache.scala 377:71]
  wire  _T_1474; // @[DCache.scala 378:79]
  wire  advance_pstore1; // @[DCache.scala 378:61]
  wire  _T_1476; // @[DCache.scala 379:34]
  reg [3:0] pstore2_way; // @[Reg.scala 11:16]
  reg [31:0] _RAND_69;
  wire [63:0] pstore1_storegen_data; // @[DCache.scala 748:27]
  reg [7:0] _T_1487; // @[Reg.scala 11:16]
  reg [31:0] _RAND_70;
  reg [7:0] _T_1493; // @[Reg.scala 11:16]
  reg [31:0] _RAND_71;
  reg [7:0] _T_1499; // @[Reg.scala 11:16]
  reg [31:0] _RAND_72;
  reg [7:0] _T_1505; // @[Reg.scala 11:16]
  reg [31:0] _RAND_73;
  reg [7:0] _T_1511; // @[Reg.scala 11:16]
  reg [31:0] _RAND_74;
  reg [7:0] _T_1517; // @[Reg.scala 11:16]
  reg [31:0] _RAND_75;
  reg [7:0] _T_1523; // @[Reg.scala 11:16]
  reg [31:0] _RAND_76;
  reg [7:0] _T_1529; // @[Reg.scala 11:16]
  reg [31:0] _RAND_77;
  wire [63:0] pstore2_storegen_data; // @[Cat.scala 30:58]
  wire [39:0] _T_1560; // @[DCache.scala 405:36]
  wire [7:0] _T_1565; // @[DCache.scala 410:47]
  wire [3:0] _T_1584; // @[Cat.scala 30:58]
  wire [3:0] _T_1587; // @[Cat.scala 30:58]
  wire [1:0] _T_1765; // @[DCache.scala 430:59]
  wire  a_source; // @[Mux.scala 31:69]
  wire [39:0] acquire_address; // @[DCache.scala 431:49]
  wire [1:0] a_size; // @[Consts.scala 19:28]
  wire [2:0] _T_1822; // @[Misc.scala 206:34]
  wire [3:0] _T_1824; // @[OneHot.scala 52:12]
  wire [2:0] _T_1826; // @[Misc.scala 206:81]
  wire  _T_1827; // @[Misc.scala 210:21]
  wire  _T_1832; // @[Misc.scala 219:38]
  wire  _T_1833; // @[Misc.scala 219:29]
  wire  _T_1835; // @[Misc.scala 219:38]
  wire  _T_1836; // @[Misc.scala 219:29]
  wire  _T_1840; // @[Misc.scala 218:27]
  wire  _T_1841; // @[Misc.scala 219:38]
  wire  _T_1842; // @[Misc.scala 219:29]
  wire  _T_1843; // @[Misc.scala 218:27]
  wire  _T_1844; // @[Misc.scala 219:38]
  wire  _T_1845; // @[Misc.scala 219:29]
  wire  _T_1846; // @[Misc.scala 218:27]
  wire  _T_1847; // @[Misc.scala 219:38]
  wire  _T_1848; // @[Misc.scala 219:29]
  wire  _T_1849; // @[Misc.scala 218:27]
  wire  _T_1850; // @[Misc.scala 219:38]
  wire  _T_1851; // @[Misc.scala 219:29]
  wire  _T_1855; // @[Misc.scala 218:27]
  wire  _T_1856; // @[Misc.scala 219:38]
  wire  _T_1857; // @[Misc.scala 219:29]
  wire  _T_1858; // @[Misc.scala 218:27]
  wire  _T_1859; // @[Misc.scala 219:38]
  wire  _T_1860; // @[Misc.scala 219:29]
  wire  _T_1861; // @[Misc.scala 218:27]
  wire  _T_1862; // @[Misc.scala 219:38]
  wire  _T_1863; // @[Misc.scala 219:29]
  wire  _T_1864; // @[Misc.scala 218:27]
  wire  _T_1865; // @[Misc.scala 219:38]
  wire  _T_1866; // @[Misc.scala 219:29]
  wire  _T_1867; // @[Misc.scala 218:27]
  wire  _T_1868; // @[Misc.scala 219:38]
  wire  _T_1869; // @[Misc.scala 219:29]
  wire  _T_1870; // @[Misc.scala 218:27]
  wire  _T_1871; // @[Misc.scala 219:38]
  wire  _T_1872; // @[Misc.scala 219:29]
  wire  _T_1873; // @[Misc.scala 218:27]
  wire  _T_1874; // @[Misc.scala 219:38]
  wire  _T_1875; // @[Misc.scala 219:29]
  wire  _T_1876; // @[Misc.scala 218:27]
  wire  _T_1877; // @[Misc.scala 219:38]
  wire  _T_1878; // @[Misc.scala 219:29]
  wire [7:0] get_mask; // @[Cat.scala 30:58]
  wire  _T_2939; // @[Mux.scala 46:19]
  wire [2:0] _T_2940_opcode; // @[Mux.scala 46:16]
  wire [2:0] _T_2940_param; // @[Mux.scala 46:16]
  wire [3:0] _T_2874_size; // @[Edges.scala 476:17 Edges.scala 479:15]
  wire [3:0] _T_2940_size; // @[Mux.scala 46:16]
  wire  _T_2940_source; // @[Mux.scala 46:16]
  wire [31:0] _T_2940_address; // @[Mux.scala 46:16]
  wire [7:0] _T_2940_mask; // @[Mux.scala 46:16]
  wire [63:0] _T_2940_data; // @[Mux.scala 46:16]
  wire  _T_2941; // @[Mux.scala 46:19]
  wire [2:0] _T_2942_opcode; // @[Mux.scala 46:16]
  wire [2:0] _T_2942_param; // @[Mux.scala 46:16]
  wire [3:0] _T_2942_size; // @[Mux.scala 46:16]
  wire  _T_2942_source; // @[Mux.scala 46:16]
  wire [31:0] _T_2942_address; // @[Mux.scala 46:16]
  wire [7:0] _T_2942_mask; // @[Mux.scala 46:16]
  wire [63:0] _T_2942_data; // @[Mux.scala 46:16]
  wire  _T_2943; // @[Mux.scala 46:19]
  wire [2:0] _T_2944_opcode; // @[Mux.scala 46:16]
  wire [2:0] _T_2944_param; // @[Mux.scala 46:16]
  wire [3:0] _T_2944_size; // @[Mux.scala 46:16]
  wire  _T_2944_source; // @[Mux.scala 46:16]
  wire [31:0] _T_2944_address; // @[Mux.scala 46:16]
  wire [7:0] _T_2944_mask; // @[Mux.scala 46:16]
  wire [63:0] _T_2944_data; // @[Mux.scala 46:16]
  wire  _T_2945; // @[Mux.scala 46:19]
  wire [2:0] _T_2946_opcode; // @[Mux.scala 46:16]
  wire [2:0] _T_2946_param; // @[Mux.scala 46:16]
  wire [3:0] _T_2946_size; // @[Mux.scala 46:16]
  wire  _T_2946_source; // @[Mux.scala 46:16]
  wire [31:0] _T_2946_address; // @[Mux.scala 46:16]
  wire [7:0] _T_2946_mask; // @[Mux.scala 46:16]
  wire [63:0] _T_2946_data; // @[Mux.scala 46:16]
  wire  _T_2947; // @[Mux.scala 46:19]
  wire [2:0] _T_2948_opcode; // @[Mux.scala 46:16]
  wire [2:0] _T_2948_param; // @[Mux.scala 46:16]
  wire [3:0] _T_2948_size; // @[Mux.scala 46:16]
  wire  _T_2948_source; // @[Mux.scala 46:16]
  wire [31:0] _T_2948_address; // @[Mux.scala 46:16]
  wire [7:0] _T_2948_mask; // @[Mux.scala 46:16]
  wire [63:0] _T_2948_data; // @[Mux.scala 46:16]
  wire  _T_2949; // @[Mux.scala 46:19]
  wire [2:0] _T_2950_opcode; // @[Mux.scala 46:16]
  wire [2:0] _T_2950_param; // @[Mux.scala 46:16]
  wire [3:0] _T_2950_size; // @[Mux.scala 46:16]
  wire  _T_2950_source; // @[Mux.scala 46:16]
  wire [31:0] _T_2950_address; // @[Mux.scala 46:16]
  wire [7:0] _T_2950_mask; // @[Mux.scala 46:16]
  wire [63:0] _T_2950_data; // @[Mux.scala 46:16]
  wire  _T_2951; // @[Mux.scala 46:19]
  wire [2:0] _T_2952_opcode; // @[Mux.scala 46:16]
  wire [2:0] _T_2952_param; // @[Mux.scala 46:16]
  wire [3:0] _T_2952_size; // @[Mux.scala 46:16]
  wire  _T_2952_source; // @[Mux.scala 46:16]
  wire [31:0] _T_2952_address; // @[Mux.scala 46:16]
  wire [7:0] _T_2952_mask; // @[Mux.scala 46:16]
  wire [63:0] _T_2952_data; // @[Mux.scala 46:16]
  wire  _T_2953; // @[Mux.scala 46:19]
  wire [2:0] _T_2954_opcode; // @[Mux.scala 46:16]
  wire [2:0] _T_2954_param; // @[Mux.scala 46:16]
  wire [3:0] _T_2954_size; // @[Mux.scala 46:16]
  wire  _T_2954_source; // @[Mux.scala 46:16]
  wire [31:0] _T_2954_address; // @[Mux.scala 46:16]
  wire [7:0] _T_2954_mask; // @[Mux.scala 46:16]
  wire [63:0] _T_2954_data; // @[Mux.scala 46:16]
  wire  _T_2955; // @[Mux.scala 46:19]
  wire [2:0] atomics_opcode; // @[Mux.scala 46:16]
  wire [2:0] atomics_param; // @[Mux.scala 46:16]
  wire [3:0] atomics_size; // @[Mux.scala 46:16]
  wire  atomics_source; // @[Mux.scala 46:16]
  wire [31:0] atomics_address; // @[Mux.scala 46:16]
  wire [7:0] atomics_mask; // @[Mux.scala 46:16]
  wire [63:0] atomics_data; // @[Mux.scala 46:16]
  wire  _T_2959; // @[DCache.scala 454:63]
  wire  tl_out_a_valid; // @[DCache.scala 454:128]
  wire [2:0] _T_3052_opcode; // @[DCache.scala 455:108]
  wire [2:0] _T_3052_param; // @[DCache.scala 455:108]
  wire [3:0] _T_3052_size; // @[DCache.scala 455:108]
  wire  _T_3052_source; // @[DCache.scala 455:108]
  wire [31:0] _T_3052_address; // @[DCache.scala 455:108]
  wire [7:0] _T_3052_mask; // @[DCache.scala 455:108]
  wire [63:0] _T_3052_data; // @[DCache.scala 455:108]
  wire [2:0] _T_3053_opcode; // @[DCache.scala 455:88]
  wire [2:0] _T_3053_param; // @[DCache.scala 455:88]
  wire [3:0] _T_3053_size; // @[DCache.scala 455:88]
  wire  _T_3053_source; // @[DCache.scala 455:88]
  wire [31:0] _T_3053_address; // @[DCache.scala 455:88]
  wire [7:0] _T_3053_mask; // @[DCache.scala 455:88]
  wire [63:0] _T_3053_data; // @[DCache.scala 455:88]
  wire [2:0] _T_2985_param; // @[Edges.scala 323:17 Edges.scala 325:15]
  wire [1:0] _T_3056; // @[OneHot.scala 52:12]
  wire  a_sel; // @[DCache.scala 458:66]
  wire  _T_3058; // @[Decoupled.scala 37:37]
  wire  _GEN_99; // @[DCache.scala 462:18]
  wire [8:0] _T_3072; // @[Edges.scala 230:28]
  wire  d_done; // @[Edges.scala 233:22]
  wire [8:0] _T_3076; // @[Edges.scala 234:25]
  wire [11:0] d_address_inc; // @[Edges.scala 269:29]
  wire  grantIsVoluntary; // @[DCache.scala 490:32]
  wire [2:0] _T_3089; // @[DCache.scala 494:97]
  wire  _T_3096; // @[DCache.scala 500:13]
  wire [1:0] _T_3099; // @[OneHot.scala 52:12]
  wire  d_sel; // @[DCache.scala 508:82]
  wire  _T_3103; // @[DCache.scala 511:17]
  wire  _T_3105; // @[DCache.scala 512:17]
  wire [31:0] dontCareBits; // @[DCache.scala 524:53]
  wire [31:0] _GEN_299; // @[DCache.scala 525:24]
  wire [31:0] _T_3110; // @[DCache.scala 525:24]
  wire  _T_3112; // @[DCache.scala 530:13]
  wire  _GEN_135; // @[DCache.scala 529:36]
  wire  _GEN_143; // @[DCache.scala 507:35]
  wire  _GEN_155; // @[DCache.scala 498:26]
  wire  _GEN_167; // @[DCache.scala 497:26]
  wire  _T_3114; // @[DCache.scala 536:36]
  wire  _T_3115; // @[DCache.scala 536:47]
  wire  tl_out__e_valid; // @[DCache.scala 544:51]
  wire  _T_3119; // @[Decoupled.scala 37:37]
  wire  _T_3121; // @[DCache.scala 538:47]
  wire  _T_3122; // @[DCache.scala 538:58]
  wire  _T_3123; // @[DCache.scala 538:26]
  wire  _T_3125; // @[DCache.scala 538:9]
  wire  _T_3127; // @[DCache.scala 543:44]
  wire [39:0] _T_3132; // @[DCache.scala 550:57]
  wire [39:0] _GEN_300; // @[DCache.scala 550:67]
  wire [39:0] _T_3133; // @[DCache.scala 550:67]
  wire  _T_3136; // @[DCache.scala 564:43]
  wire [3:0] _T_3195; // @[Cat.scala 30:58]
  wire  _T_3204; // @[Mux.scala 46:19]
  wire [1:0] _T_3205; // @[Mux.scala 46:16]
  wire  _T_3206; // @[Mux.scala 46:19]
  wire [1:0] _T_3207; // @[Mux.scala 46:16]
  wire  _T_3208; // @[Mux.scala 46:19]
  wire [1:0] _T_3209; // @[Mux.scala 46:16]
  wire  _T_3210; // @[Mux.scala 46:19]
  wire [1:0] _T_3211; // @[Mux.scala 46:16]
  wire  _GEN_170; // @[DCache.scala 577:27]
  wire  _GEN_171; // @[DCache.scala 577:27]
  wire  _GEN_172; // @[DCache.scala 577:27]
  wire  _T_3227; // @[DCache.scala 588:61]
  wire  _T_3228; // @[DCache.scala 588:44]
  wire [39:0] _T_3237; // @[Cat.scala 30:58]
  wire [8:0] _T_3250; // @[Edges.scala 230:28]
  wire  c_first; // @[Edges.scala 231:25]
  wire [8:0] c_count; // @[Edges.scala 234:25]
  wire  releaseRejected; // @[DCache.scala 598:40]
  reg  s1_release_data_valid; // @[DCache.scala 599:34]
  reg [31:0] _RAND_78;
  wire [9:0] _T_3261; // @[Cat.scala 30:58]
  wire [1:0] _T_3262; // @[Cat.scala 30:58]
  wire [1:0] _GEN_301; // @[DCache.scala 601:101]
  wire [1:0] _T_3264; // @[DCache.scala 601:101]
  wire [1:0] _T_3265; // @[DCache.scala 601:52]
  wire [9:0] _GEN_302; // @[DCache.scala 601:47]
  wire [9:0] releaseDataBeat; // @[DCache.scala 601:47]
  wire  _T_3291; // @[DCache.scala 615:24]
  wire  _T_3292; // @[DCache.scala 616:25]
  wire  _T_3297; // @[DCache.scala 616:13]
  wire [25:0] _T_3300; // @[Cat.scala 30:58]
  wire [31:0] res_2_address; // @[DCache.scala 618:96]
  wire [2:0] _GEN_180; // @[DCache.scala 615:44]
  wire [2:0] _T_3305; // @[DCache.scala 629:29]
  wire [2:0] _T_3307; // @[DCache.scala 633:29]
  wire [2:0] _GEN_191; // @[DCache.scala 626:45]
  wire [2:0] _GEN_197; // @[DCache.scala 626:45]
  wire [2:0] _GEN_199; // @[DCache.scala 624:36]
  wire [2:0] _GEN_202; // @[DCache.scala 624:36]
  wire [2:0] _GEN_220; // @[DCache.scala 620:21]
  wire [2:0] _GEN_223; // @[DCache.scala 620:21]
  wire  _T_3308; // @[DCache.scala 637:25]
  wire [39:0] _T_3311; // @[Cat.scala 30:58]
  wire [2:0] _GEN_230; // @[DCache.scala 641:37]
  wire  _GEN_231; // @[DCache.scala 641:37]
  wire [2:0] _GEN_235; // @[DCache.scala 637:44]
  wire [2:0] _GEN_237; // @[DCache.scala 648:26]
  wire [2:0] _GEN_239; // @[DCache.scala 646:47]
  wire [2:0] _GEN_243; // @[DCache.scala 650:48]
  wire [2:0] _GEN_252; // @[DCache.scala 655:48]
  wire  _T_3340; // @[DCache.scala 668:29]
  wire  _GEN_260; // @[DCache.scala 668:41]
  wire [1:0] newCoh_state; // @[DCache.scala 659:81]
  wire  _T_3342; // @[DCache.scala 676:60]
  wire [11:0] _T_3345; // @[DCache.scala 679:55]
  wire [5:0] _T_3347; // @[DCache.scala 679:117]
  wire [11:0] _GEN_304; // @[DCache.scala 679:72]
  wire  _T_3352; // @[package.scala 14:47]
  wire  _T_3362; // @[Decoupled.scala 37:37]
  wire  _T_3367; // @[DCache.scala 701:57]
  wire  _T_3368; // @[DCache.scala 701:94]
  wire  _T_3370; // @[DCache.scala 701:115]
  reg  _T_3374; // @[DCache.scala 705:32]
  reg [31:0] _RAND_79;
  reg  _T_3376_pf_ld; // @[Reg.scala 11:16]
  reg [31:0] _RAND_80;
  reg  _T_3376_pf_st; // @[Reg.scala 11:16]
  reg [31:0] _RAND_81;
  reg  _T_3376_ae_ld; // @[Reg.scala 11:16]
  reg [31:0] _RAND_82;
  reg  _T_3376_ae_st; // @[Reg.scala 11:16]
  reg [31:0] _RAND_83;
  reg  _T_3376_ma_ld; // @[Reg.scala 11:16]
  reg [31:0] _RAND_84;
  reg  _T_3376_ma_st; // @[Reg.scala 11:16]
  reg [31:0] _RAND_85;
  reg  doUncachedResp; // @[DCache.scala 720:27]
  reg [31:0] _RAND_86;
  wire  _T_3403; // @[DCache.scala 723:11]
  wire [31:0] _T_3412; // @[AMOALU.scala 39:24]
  wire  _T_3415; // @[AMOALU.scala 42:26]
  wire  _T_3418; // @[AMOALU.scala 42:76]
  wire [31:0] _T_3420; // @[Bitwise.scala 72:12]
  wire [31:0] _T_3422; // @[AMOALU.scala 42:20]
  wire [63:0] _T_3423; // @[Cat.scala 30:58]
  wire [15:0] _T_3427; // @[AMOALU.scala 39:24]
  wire  _T_3430; // @[AMOALU.scala 42:26]
  wire  _T_3433; // @[AMOALU.scala 42:76]
  wire [47:0] _T_3435; // @[Bitwise.scala 72:12]
  wire [47:0] _T_3437; // @[AMOALU.scala 42:20]
  wire [63:0] _T_3438; // @[Cat.scala 30:58]
  wire [7:0] _T_3442; // @[AMOALU.scala 39:24]
  wire [7:0] _T_3444; // @[AMOALU.scala 41:23]
  wire  _T_3445; // @[AMOALU.scala 42:26]
  wire  _T_3446; // @[AMOALU.scala 42:38]
  wire  _T_3448; // @[AMOALU.scala 42:76]
  wire [55:0] _T_3450; // @[Bitwise.scala 72:12]
  wire [55:0] _T_3452; // @[AMOALU.scala 42:20]
  wire [63:0] _T_3453; // @[Cat.scala 30:58]
  wire [63:0] _GEN_305; // @[DCache.scala 735:41]
  reg  resetting; // @[DCache.scala 757:26]
  reg [31:0] _RAND_87;
  reg  _T_3473; // @[DCache.scala 759:18]
  reg [31:0] _RAND_88;
  wire  _GEN_290; // @[DCache.scala 759:27]
  reg  flushed; // @[DCache.scala 760:20]
  reg [31:0] _RAND_89;
  reg  flushing; // @[DCache.scala 761:21]
  reg [31:0] _RAND_90;
  reg [7:0] flushCounter; // @[DCache.scala 762:25]
  reg [31:0] _RAND_91;
  wire [8:0] flushCounterNext; // @[DCache.scala 763:39]
  wire  flushDone; // @[DCache.scala 764:57]
  wire  _T_3478; // @[DCache.scala 766:39]
  wire  _T_3479; // @[DCache.scala 766:25]
  wire  _T_3487; // @[DCache.scala 769:56]
  wire  _T_3494; // @[Decoupled.scala 37:37]
  wire  _T_3496; // @[DCache.scala 774:45]
  wire  _T_3498; // @[DCache.scala 774:64]
  wire  _T_3500; // @[DCache.scala 774:95]
  wire [11:0] _T_3505; // @[DCache.scala 778:98]
  wire [8:0] _GEN_295; // @[DCache.scala 805:20]
  wire  _T_3516; // @[DCache.scala 815:31]
  wire  _T_3517; // @[DCache.scala 816:26]
  wire  _T_3518; // @[DCache.scala 817:14]
  wire  _T_3519; // @[DCache.scala 817:26]
  wire  _T_3520; // @[DCache.scala 818:14]
  wire  _T_3521; // @[DCache.scala 818:35]
  wire  _T_3522; // @[DCache.scala 819:18]
  wire  _T_3524; // @[DCache.scala 819:35]
  wire  _T_3525; // @[DCache.scala 820:31]
  wire  _T_3529; // @[DCache.scala 821:46]
  wire  _T_3530; // @[DCache.scala 822:23]
  wire  _T_3532; // @[DCache.scala 823:23]
  wire  _T_3534; // @[DCache.scala 823:54]
  wire  _GEN_308; // @[DCache.scala 500:13]
  wire  _GEN_311; // @[DCache.scala 512:17]
  wire  _GEN_312; // @[DCache.scala 512:17]
  wire  _GEN_313; // @[DCache.scala 512:17]
  wire  _GEN_321; // @[DCache.scala 530:13]
  wire  _GEN_322; // @[DCache.scala 530:13]
  reg [19:0] DCache_state; // @[Register tracking DCache state]
  reg [31:0] _RAND_92;
  reg  DCache_cov [0:1048575]; // @[Coverage map for DCache]
  reg [31:0] _RAND_93;
  wire  DCache_cov_read_data; // @[Coverage map for DCache]
  wire [19:0] DCache_cov_read_addr; // @[Coverage map for DCache]
  wire  DCache_cov_write_data; // @[Coverage map for DCache]
  wire [19:0] DCache_cov_write_addr; // @[Coverage map for DCache]
  wire  DCache_cov_write_mask; // @[Coverage map for DCache]
  wire  DCache_cov_write_en; // @[Coverage map for DCache]
  reg [29:0] DCache_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_94;
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  mux_cond_4;
  wire  mux_cond_5;
  wire [18:0] pstore1_held_shl;
  wire [19:0] pstore1_held_pad;
  wire [15:0] s2_valid_pre_xcpt_shl;
  wire [19:0] s2_valid_pre_xcpt_pad;
  wire [7:0] s2_release_data_valid_shl;
  wire [19:0] s2_release_data_valid_pad;
  wire [15:0] s2_flush_valid_pre_tag_ecc_shl;
  wire [19:0] s2_flush_valid_pre_tag_ecc_pad;
  wire [14:0] s2_hit_way_shl;
  wire [19:0] s2_hit_way_pad;
  wire [4:0] _T_1060_shl;
  wire [19:0] _T_1060_pad;
  wire [12:0] s2_hit_state_state_shl;
  wire [19:0] s2_hit_state_state_pad;
  wire [18:0] pstore2_valid_shl;
  wire [19:0] pstore2_valid_pad;
  wire [15:0] uncachedInFlight_0_shl;
  wire [19:0] uncachedInFlight_0_pad;
  wire [6:0] s2_probe_shl;
  wire [19:0] s2_probe_pad;
  wire [12:0] resetting_shl;
  wire [19:0] resetting_pad;
  wire [4:0] s2_probe_way_shl;
  wire [19:0] s2_probe_way_pad;
  wire [12:0] s1_valid_shl;
  wire [19:0] s1_valid_pad;
  wire [18:0] grantInProgress_shl;
  wire [19:0] grantInProgress_pad;
  wire [10:0] s2_req_typ_shl;
  wire [19:0] s2_req_typ_pad;
  wire [1:0] s2_probe_state_state_shl;
  wire [19:0] s2_probe_state_state_pad;
  wire [3:0] cached_grant_wait_shl;
  wire [19:0] cached_grant_wait_pad;
  wire [12:0] flushed_shl;
  wire [19:0] flushed_pad;
  wire [5:0] release_ack_wait_shl;
  wire [19:0] release_ack_wait_pad;
  wire [15:0] s2_uncached_shl;
  wire [19:0] s2_uncached_pad;
  wire [19:0] release_state_shl;
  wire [19:0] release_state_pad;
  wire [16:0] s1_flush_valid_shl;
  wire [19:0] s1_flush_valid_pad;
  wire [4:0] blockUncachedGrant_shl;
  wire [19:0] blockUncachedGrant_pad;
  wire [1:0] _T_1068_state_shl;
  wire [19:0] _T_1068_state_pad;
  wire [1:0] _T_738_shl;
  wire [19:0] _T_738_pad;
  wire [15:0] probe_bits_param_shl;
  wire [19:0] probe_bits_param_pad;
  wire [4:0] s1_probe_shl;
  wire [19:0] s1_probe_pad;
  wire [6:0] pstore1_rmw_shl;
  wire [19:0] pstore1_rmw_pad;
  wire [16:0] s1_req_typ_shl;
  wire [19:0] s1_req_typ_pad;
  wire [11:0] mux_cond_0_shl;
  wire [19:0] mux_cond_0_pad;
  wire [10:0] mux_cond_1_shl;
  wire [19:0] mux_cond_1_pad;
  wire [1:0] mux_cond_2_shl;
  wire [19:0] mux_cond_2_pad;
  wire [12:0] mux_cond_3_shl;
  wire [19:0] mux_cond_3_pad;
  wire [17:0] mux_cond_4_shl;
  wire [19:0] mux_cond_4_pad;
  wire [2:0] mux_cond_5_shl;
  wire [19:0] mux_cond_5_pad;
  wire [19:0] DCache_xor15;
  wire [19:0] DCache_xor16;
  wire [19:0] DCache_xor7;
  wire [19:0] DCache_xor17;
  wire [19:0] DCache_xor18;
  wire [19:0] DCache_xor8;
  wire [19:0] DCache_xor3;
  wire [19:0] DCache_xor19;
  wire [19:0] DCache_xor20;
  wire [19:0] DCache_xor9;
  wire [19:0] DCache_xor21;
  wire [19:0] DCache_xor46;
  wire [19:0] DCache_xor22;
  wire [19:0] DCache_xor10;
  wire [19:0] DCache_xor4;
  wire [19:0] DCache_xor1;
  wire [19:0] DCache_xor23;
  wire [19:0] DCache_xor24;
  wire [19:0] DCache_xor11;
  wire [19:0] DCache_xor25;
  wire [19:0] DCache_xor54;
  wire [19:0] DCache_xor26;
  wire [19:0] DCache_xor12;
  wire [19:0] DCache_xor5;
  wire [19:0] DCache_xor27;
  wire [19:0] DCache_xor28;
  wire [19:0] DCache_xor13;
  wire [19:0] DCache_xor29;
  wire [19:0] DCache_xor62;
  wire [19:0] DCache_xor30;
  wire [19:0] DCache_xor14;
  wire [19:0] DCache_xor6;
  wire [19:0] DCache_xor2;
  wire [19:0] DCache_xor0;
  wire [29:0] dataArb_sum;
  wire [29:0] amoalu_sum;
  wire [29:0] data_sum;
  wire [29:0] metaArb_sum;
  wire [29:0] tlb_sum;
  wire  stopEn0;
  wire  stopEn1;
  wire  stopEn2;
  wire  stopEn3;
  wire  stopEn4;
  wire  stopEn5;
  wire  stopEn6;
  wire  stopEn7;
  wire  stopEn8;
  wire  dataArb_metaAssert_wire;
  wire  metaArb_metaAssert_wire;
  wire  tlb_metaAssert_wire;
  wire  data_metaAssert_wire;
  wire  amoalu_metaAssert_wire;
  wire  DCache_or8;
  wire  DCache_or3;
  wire  DCache_or9;
  wire  DCache_or10;
  wire  DCache_or4;
  wire  DCache_or1;
  wire  DCache_or12;
  wire  DCache_or5;
  wire  DCache_or13;
  wire  DCache_or14;
  wire  DCache_or6;
  wire  DCache_or2;
  wire  DCache_or0;
  Arbiter metaArb ( // @[DCache.scala 98:23]
    .io_in_0_valid(metaArb_io_in_0_valid),
    .io_in_0_bits_addr(metaArb_io_in_0_bits_addr),
    .io_in_0_bits_idx(metaArb_io_in_0_bits_idx),
    .io_in_0_bits_data(metaArb_io_in_0_bits_data),
    .io_in_2_valid(metaArb_io_in_2_valid),
    .io_in_2_bits_addr(metaArb_io_in_2_bits_addr),
    .io_in_2_bits_idx(metaArb_io_in_2_bits_idx),
    .io_in_2_bits_way_en(metaArb_io_in_2_bits_way_en),
    .io_in_2_bits_data(metaArb_io_in_2_bits_data),
    .io_in_3_valid(metaArb_io_in_3_valid),
    .io_in_3_bits_addr(metaArb_io_in_3_bits_addr),
    .io_in_3_bits_idx(metaArb_io_in_3_bits_idx),
    .io_in_3_bits_way_en(metaArb_io_in_3_bits_way_en),
    .io_in_3_bits_data(metaArb_io_in_3_bits_data),
    .io_in_4_ready(metaArb_io_in_4_ready),
    .io_in_4_valid(metaArb_io_in_4_valid),
    .io_in_4_bits_addr(metaArb_io_in_4_bits_addr),
    .io_in_4_bits_idx(metaArb_io_in_4_bits_idx),
    .io_in_4_bits_way_en(metaArb_io_in_4_bits_way_en),
    .io_in_4_bits_data(metaArb_io_in_4_bits_data),
    .io_in_5_ready(metaArb_io_in_5_ready),
    .io_in_5_valid(metaArb_io_in_5_valid),
    .io_in_5_bits_addr(metaArb_io_in_5_bits_addr),
    .io_in_5_bits_idx(metaArb_io_in_5_bits_idx),
    .io_in_5_bits_way_en(metaArb_io_in_5_bits_way_en),
    .io_in_5_bits_data(metaArb_io_in_5_bits_data),
    .io_in_6_ready(metaArb_io_in_6_ready),
    .io_in_6_valid(metaArb_io_in_6_valid),
    .io_in_6_bits_addr(metaArb_io_in_6_bits_addr),
    .io_in_6_bits_idx(metaArb_io_in_6_bits_idx),
    .io_in_6_bits_way_en(metaArb_io_in_6_bits_way_en),
    .io_in_6_bits_data(metaArb_io_in_6_bits_data),
    .io_in_7_ready(metaArb_io_in_7_ready),
    .io_in_7_valid(metaArb_io_in_7_valid),
    .io_in_7_bits_addr(metaArb_io_in_7_bits_addr),
    .io_in_7_bits_idx(metaArb_io_in_7_bits_idx),
    .io_in_7_bits_way_en(metaArb_io_in_7_bits_way_en),
    .io_in_7_bits_data(metaArb_io_in_7_bits_data),
    .io_out_ready(metaArb_io_out_ready),
    .io_out_valid(metaArb_io_out_valid),
    .io_out_bits_write(metaArb_io_out_bits_write),
    .io_out_bits_addr(metaArb_io_out_bits_addr),
    .io_out_bits_idx(metaArb_io_out_bits_idx),
    .io_out_bits_way_en(metaArb_io_out_bits_way_en),
    .io_out_bits_data(metaArb_io_out_bits_data),
    .io_covSum(metaArb_io_covSum),
    .metaAssert(metaArb_metaAssert)
  );
  DCacheDataArray data ( // @[DCache.scala 108:20]
    .clock(data_clock),
    .io_req_valid(data_io_req_valid),
    .io_req_bits_addr(data_io_req_bits_addr),
    .io_req_bits_write(data_io_req_bits_write),
    .io_req_bits_wdata(data_io_req_bits_wdata),
    .io_req_bits_eccMask(data_io_req_bits_eccMask),
    .io_req_bits_way_en(data_io_req_bits_way_en),
    .io_resp_0(data_io_resp_0),
    .io_resp_1(data_io_resp_1),
    .io_resp_2(data_io_resp_2),
    .io_resp_3(data_io_resp_3),
    .io_covSum(data_io_covSum),
    .metaAssert(data_metaAssert),
    .metaReset(data_metaReset)
  );
  Arbiter_1 dataArb ( // @[DCache.scala 109:23]
    .io_in_0_valid(dataArb_io_in_0_valid),
    .io_in_0_bits_addr(dataArb_io_in_0_bits_addr),
    .io_in_0_bits_write(dataArb_io_in_0_bits_write),
    .io_in_0_bits_wdata(dataArb_io_in_0_bits_wdata),
    .io_in_0_bits_eccMask(dataArb_io_in_0_bits_eccMask),
    .io_in_0_bits_way_en(dataArb_io_in_0_bits_way_en),
    .io_in_1_ready(dataArb_io_in_1_ready),
    .io_in_1_valid(dataArb_io_in_1_valid),
    .io_in_1_bits_addr(dataArb_io_in_1_bits_addr),
    .io_in_1_bits_write(dataArb_io_in_1_bits_write),
    .io_in_1_bits_wdata(dataArb_io_in_1_bits_wdata),
    .io_in_1_bits_eccMask(dataArb_io_in_1_bits_eccMask),
    .io_in_1_bits_way_en(dataArb_io_in_1_bits_way_en),
    .io_in_2_ready(dataArb_io_in_2_ready),
    .io_in_2_valid(dataArb_io_in_2_valid),
    .io_in_2_bits_addr(dataArb_io_in_2_bits_addr),
    .io_in_2_bits_wdata(dataArb_io_in_2_bits_wdata),
    .io_in_2_bits_eccMask(dataArb_io_in_2_bits_eccMask),
    .io_in_3_ready(dataArb_io_in_3_ready),
    .io_in_3_valid(dataArb_io_in_3_valid),
    .io_in_3_bits_addr(dataArb_io_in_3_bits_addr),
    .io_in_3_bits_wdata(dataArb_io_in_3_bits_wdata),
    .io_in_3_bits_eccMask(dataArb_io_in_3_bits_eccMask),
    .io_out_valid(dataArb_io_out_valid),
    .io_out_bits_addr(dataArb_io_out_bits_addr),
    .io_out_bits_write(dataArb_io_out_bits_write),
    .io_out_bits_wdata(dataArb_io_out_bits_wdata),
    .io_out_bits_eccMask(dataArb_io_out_bits_eccMask),
    .io_out_bits_way_en(dataArb_io_out_bits_way_en),
    .io_covSum(dataArb_io_covSum),
    .metaAssert(dataArb_metaAssert)
  );
  TLB tlb ( // @[DCache.scala 184:19]
    .clock(tlb_clock),
    .reset(tlb_reset),
    .io_req_ready(tlb_io_req_ready),
    .io_req_valid(tlb_io_req_valid),
    .io_req_bits_vaddr(tlb_io_req_bits_vaddr),
    .io_req_bits_passthrough(tlb_io_req_bits_passthrough),
    .io_req_bits_size(tlb_io_req_bits_size),
    .io_req_bits_cmd(tlb_io_req_bits_cmd),
    .io_resp_miss(tlb_io_resp_miss),
    .io_resp_paddr(tlb_io_resp_paddr),
    .io_resp_pf_ld(tlb_io_resp_pf_ld),
    .io_resp_pf_st(tlb_io_resp_pf_st),
    .io_resp_ae_ld(tlb_io_resp_ae_ld),
    .io_resp_ae_st(tlb_io_resp_ae_st),
    .io_resp_ma_ld(tlb_io_resp_ma_ld),
    .io_resp_ma_st(tlb_io_resp_ma_st),
    .io_resp_cacheable(tlb_io_resp_cacheable),
    .io_sfence_valid(tlb_io_sfence_valid),
    .io_sfence_bits_rs1(tlb_io_sfence_bits_rs1),
    .io_sfence_bits_rs2(tlb_io_sfence_bits_rs2),
    .io_sfence_bits_addr(tlb_io_sfence_bits_addr),
    .io_ptw_req_ready(tlb_io_ptw_req_ready),
    .io_ptw_req_valid(tlb_io_ptw_req_valid),
    .io_ptw_req_bits_valid(tlb_io_ptw_req_bits_valid),
    .io_ptw_req_bits_bits_addr(tlb_io_ptw_req_bits_bits_addr),
    .io_ptw_resp_valid(tlb_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae(tlb_io_ptw_resp_bits_ae),
    .io_ptw_resp_bits_pte_ppn(tlb_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d(tlb_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(tlb_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(tlb_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(tlb_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(tlb_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(tlb_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(tlb_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(tlb_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(tlb_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous(tlb_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(tlb_io_ptw_ptbr_mode),
    .io_ptw_status_dprv(tlb_io_ptw_status_dprv),
    .io_ptw_status_mxr(tlb_io_ptw_status_mxr),
    .io_ptw_status_sum(tlb_io_ptw_status_sum),
    .io_ptw_pmp_0_cfg_l(tlb_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a(tlb_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(tlb_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(tlb_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(tlb_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(tlb_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(tlb_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(tlb_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a(tlb_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(tlb_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(tlb_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(tlb_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(tlb_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(tlb_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(tlb_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a(tlb_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(tlb_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(tlb_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(tlb_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(tlb_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(tlb_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(tlb_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a(tlb_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(tlb_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(tlb_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(tlb_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(tlb_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(tlb_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(tlb_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a(tlb_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(tlb_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(tlb_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(tlb_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(tlb_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(tlb_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(tlb_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a(tlb_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(tlb_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(tlb_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(tlb_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(tlb_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(tlb_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(tlb_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a(tlb_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(tlb_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(tlb_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(tlb_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(tlb_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(tlb_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(tlb_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a(tlb_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(tlb_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(tlb_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(tlb_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(tlb_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(tlb_io_ptw_pmp_7_mask),
    .io_ptw_vpoffset_bits_value(tlb_io_ptw_vpoffset_bits_value),
    .io_covSum(tlb_io_covSum),
    .metaAssert(tlb_metaAssert),
    .metaReset(tlb_metaReset)
  );
  AMOALU amoalu ( // @[DCache.scala 743:24]
    .io_mask(amoalu_io_mask),
    .io_cmd(amoalu_io_cmd),
    .io_lhs(amoalu_io_lhs),
    .io_rhs(amoalu_io_rhs),
    .io_out(amoalu_io_out),
    .io_covSum(amoalu_io_covSum),
    .metaAssert(amoalu_metaAssert)
  );
  assign tag_array_0_s1_meta_addr = tag_array_0_s1_meta_addr_pipe_0;
  assign tag_array_0_s1_meta_data = tag_array_0[tag_array_0_s1_meta_addr]; // @[DescribedSRAM.scala 23:21]
  assign tag_array_0__T_567_data = metaArb_io_out_bits_data;
  assign tag_array_0__T_567_addr = metaArb_io_out_bits_idx;
  assign tag_array_0__T_567_mask = metaArb_io_out_bits_way_en[0];
  assign tag_array_0__T_567_en = metaArb_io_out_valid & metaArb_io_out_bits_write;
  assign tag_array_1_s1_meta_addr = tag_array_1_s1_meta_addr_pipe_0;
  assign tag_array_1_s1_meta_data = tag_array_1[tag_array_1_s1_meta_addr]; // @[DescribedSRAM.scala 23:21]
  assign tag_array_1__T_567_data = metaArb_io_out_bits_data;
  assign tag_array_1__T_567_addr = metaArb_io_out_bits_idx;
  assign tag_array_1__T_567_mask = metaArb_io_out_bits_way_en[1];
  assign tag_array_1__T_567_en = metaArb_io_out_valid & metaArb_io_out_bits_write;
  assign tag_array_2_s1_meta_addr = tag_array_2_s1_meta_addr_pipe_0;
  assign tag_array_2_s1_meta_data = tag_array_2[tag_array_2_s1_meta_addr]; // @[DescribedSRAM.scala 23:21]
  assign tag_array_2__T_567_data = metaArb_io_out_bits_data;
  assign tag_array_2__T_567_addr = metaArb_io_out_bits_idx;
  assign tag_array_2__T_567_mask = metaArb_io_out_bits_way_en[2];
  assign tag_array_2__T_567_en = metaArb_io_out_valid & metaArb_io_out_bits_write;
  assign tag_array_3_s1_meta_addr = tag_array_3_s1_meta_addr_pipe_0;
  assign tag_array_3_s1_meta_data = tag_array_3[tag_array_3_s1_meta_addr]; // @[DescribedSRAM.scala 23:21]
  assign tag_array_3__T_567_data = metaArb_io_out_bits_data;
  assign tag_array_3__T_567_addr = metaArb_io_out_bits_idx;
  assign tag_array_3__T_567_mask = metaArb_io_out_bits_way_en[3];
  assign tag_array_3__T_567_en = metaArb_io_out_valid & metaArb_io_out_bits_write;
  assign _T_251 = lfsr[0] ^ lfsr[2]; // @[LFSR.scala 23:43]
  assign _T_253 = _T_251 ^ lfsr[3]; // @[LFSR.scala 23:51]
  assign _T_255 = _T_253 ^ lfsr[5]; // @[LFSR.scala 23:59]
  assign _T_257 = {_T_255,lfsr[15:1]}; // @[Cat.scala 30:58]
  assign grantIsUncachedData = auto_out_d_bits_opcode == 3'h1; // @[package.scala 14:47]
  assign _T_3218 = blockUncachedGrant | s1_valid; // @[DCache.scala 574:52]
  assign _T_3219 = grantIsUncachedData & _T_3218; // @[DCache.scala 574:29]
  assign grantIsRefill = auto_out_d_bits_opcode == 3'h5; // @[DCache.scala 491:29]
  assign _T_3130 = grantIsRefill & ~dataArb_io_in_1_ready; // @[DCache.scala 544:23]
  assign _T_3082 = auto_out_d_bits_opcode == 3'h4; // @[package.scala 14:47]
  assign grantIsCached = _T_3082 | grantIsRefill; // @[package.scala 14:62]
  assign d_first = _T_3069 == 9'h0; // @[Edges.scala 231:25]
  assign _T_3091 = ~d_first | auto_out_e_ready; // @[DCache.scala 496:50]
  assign _T_3093 = grantIsCached ? _T_3091 : 1'h1; // @[DCache.scala 496:24]
  assign _GEN_169 = _T_3130 ? 1'h0 : _T_3093; // @[DCache.scala 544:51]
  assign tl_out__d_ready = _T_3219 ? 1'h0 : _GEN_169; // @[DCache.scala 574:66]
  assign _T_3094 = tl_out__d_ready & auto_out_d_valid; // @[Decoupled.scala 37:37]
  assign _T_3073 = _T_3069 == 9'h1; // @[Edges.scala 232:25]
  assign _T_3062 = 27'hfff << auto_out_d_bits_size; // @[package.scala 185:77]
  assign _T_3065 = ~_T_3062[11:3]; // @[Edges.scala 220:59]
  assign _T_3067 = auto_out_d_bits_opcode[0] ? _T_3065 : 9'h0; // @[Edges.scala 221:14]
  assign _T_3074 = _T_3067 == 9'h0; // @[Edges.scala 232:47]
  assign d_last = _T_3073 | _T_3074; // @[Edges.scala 232:37]
  assign _GEN_147 = grantIsCached & d_last; // @[DCache.scala 498:26]
  assign _GEN_159 = _T_3094 & _GEN_147; // @[DCache.scala 497:26]
  assign _T_270 = dataArb_io_out_bits_wdata; // @[DCache.scala 112:65]
  assign _T_281 = {_T_270[31:24],_T_270[23:16],_T_270[15:8],_T_270[7:0]}; // @[Cat.scala 30:58]
  assign _T_284 = {_T_270[63:56],_T_270[55:48],_T_270[47:40],_T_270[39:32]}; // @[Cat.scala 30:58]
  assign _T_288 = io_cpu_req_ready & io_cpu_req_valid; // @[Decoupled.scala 37:37]
  assign _T_734 = s1_probe | s2_probe; // @[DCache.scala 233:34]
  assign _T_735 = release_state != 3'h0; // @[DCache.scala 233:63]
  assign releaseInFlight = _T_734 | _T_735; // @[DCache.scala 233:46]
  assign _T_3223 = releaseInFlight | grantInProgress; // @[DCache.scala 587:37]
  assign _T_3224 = blockProbeAfterGrantCount > 3'h0; // @[DCache.scala 587:85]
  assign _T_3225 = _T_3223 | _T_3224; // @[DCache.scala 587:56]
  assign lrscValid = lrscCount > 7'h3; // @[DCache.scala 328:29]
  assign block_probe = _T_3225 | lrscValid; // @[DCache.scala 587:89]
  assign _T_3230 = metaArb_io_in_6_ready & ~block_probe; // @[DCache.scala 589:44]
  assign _T_3232 = _T_3230 & ~s1_valid; // @[DCache.scala 589:60]
  assign _T_730 = {io_cpu_s2_xcpt_ma_ld,io_cpu_s2_xcpt_ma_st,io_cpu_s2_xcpt_pf_ld,io_cpu_s2_xcpt_pf_st,io_cpu_s2_xcpt_ae_ld,io_cpu_s2_xcpt_ae_st}; // @[DCache.scala 231:55]
  assign _T_731 = _T_730 != 6'h0; // @[DCache.scala 231:62]
  assign s2_valid = s2_valid_pre_xcpt & ~_T_731; // @[DCache.scala 231:36]
  assign tl_out__b_ready = _T_3232 & ~s2_valid; // @[DCache.scala 589:73]
  assign _T_290 = tl_out__b_ready & auto_out_b_valid; // @[Decoupled.scala 37:37]
  assign s1_valid_masked = s1_valid & ~io_cpu_s1_kill; // @[DCache.scala 135:34]
  assign _T_1069 = {probe_bits_param,s2_probe_state_state}; // @[Cat.scala 30:58]
  assign _T_1126 = 4'h3 == _T_1069; // @[Misc.scala 58:20]
  assign _T_1122 = 4'h2 == _T_1069; // @[Misc.scala 58:20]
  assign _T_1118 = 4'h1 == _T_1069; // @[Misc.scala 58:20]
  assign _T_1114 = 4'h0 == _T_1069; // @[Misc.scala 58:20]
  assign _T_1110 = 4'h7 == _T_1069; // @[Misc.scala 58:20]
  assign _T_1106 = 4'h6 == _T_1069; // @[Misc.scala 58:20]
  assign _T_1102 = 4'h5 == _T_1069; // @[Misc.scala 58:20]
  assign _T_1098 = 4'h4 == _T_1069; // @[Misc.scala 58:20]
  assign _T_1094 = 4'hb == _T_1069; // @[Misc.scala 58:20]
  assign _T_1090 = 4'ha == _T_1069; // @[Misc.scala 58:20]
  assign _T_1086 = 4'h9 == _T_1069; // @[Misc.scala 58:20]
  assign _T_1082 = 4'h8 == _T_1069; // @[Misc.scala 58:20]
  assign _T_1099 = _T_1098 ? 1'h0 : _T_1094; // @[Misc.scala 40:9]
  assign _T_1103 = _T_1102 ? 1'h0 : _T_1099; // @[Misc.scala 40:9]
  assign _T_1107 = _T_1106 ? 1'h0 : _T_1103; // @[Misc.scala 40:9]
  assign _T_1111 = _T_1110 | _T_1107; // @[Misc.scala 40:9]
  assign _T_1115 = _T_1114 ? 1'h0 : _T_1111; // @[Misc.scala 40:9]
  assign _T_1119 = _T_1118 ? 1'h0 : _T_1115; // @[Misc.scala 40:9]
  assign _T_1123 = _T_1122 ? 1'h0 : _T_1119; // @[Misc.scala 40:9]
  assign s2_prb_ack_data = _T_1126 | _T_1123; // @[Misc.scala 40:9]
  assign _T_3304 = s2_probe_state_state > 2'h0; // @[Metadata.scala 50:45]
  assign _T_3251 = _T_3247 == 9'h1; // @[Edges.scala 232:25]
  assign _T_3315 = release_state == 3'h1; // @[package.scala 14:47]
  assign _T_3316 = release_state == 3'h6; // @[package.scala 14:47]
  assign _T_3317 = _T_3315 | _T_3316; // @[package.scala 14:62]
  assign _T_3314 = release_state == 3'h2; // @[DCache.scala 655:25]
  assign _T_3313 = release_state == 3'h3; // @[DCache.scala 650:25]
  assign _GEN_251 = _T_3314 ? 3'h5 : 3'h4; // @[DCache.scala 655:48]
  assign tl_out__c_bits_opcode = _T_3317 ? 3'h7 : _GEN_251; // @[DCache.scala 659:81]
  assign tl_out__c_bits_size = _T_3317 ? 4'h6 : probe_bits_size; // @[DCache.scala 659:81]
  assign _T_3240 = 27'hfff << tl_out__c_bits_size; // @[package.scala 185:77]
  assign _T_3243 = ~_T_3240[11:3]; // @[Edges.scala 220:59]
  assign _T_3245 = tl_out__c_bits_opcode[0] ? _T_3243 : 9'h0; // @[Edges.scala 221:14]
  assign _T_3252 = _T_3245 == 9'h0; // @[Edges.scala 232:47]
  assign c_last = _T_3251 | _T_3252; // @[Edges.scala 232:37]
  assign _T_3312 = release_state == 3'h5; // @[DCache.scala 646:25]
  assign _GEN_200 = s2_prb_ack_data ? s2_release_data_valid : 1'h1; // @[DCache.scala 624:36]
  assign _GEN_221 = s2_probe ? _GEN_200 : s2_release_data_valid; // @[DCache.scala 620:21]
  assign _GEN_238 = _T_3312 | _GEN_221; // @[DCache.scala 646:47]
  assign tl_out__c_valid = _T_3313 | _GEN_238; // @[DCache.scala 650:48]
  assign _T_3238 = auto_out_c_ready & tl_out__c_valid; // @[Decoupled.scala 37:37]
  assign releaseDone = c_last & _T_3238; // @[Edges.scala 233:22]
  assign _GEN_198 = _T_3304 | ~releaseDone; // @[DCache.scala 626:45]
  assign probeNack = s2_prb_ack_data | _GEN_198; // @[DCache.scala 624:36]
  assign _T_302 = s1_req_cmd == 5'h0; // @[Consts.scala 93:31]
  assign _T_303 = s1_req_cmd == 5'h6; // @[Consts.scala 93:48]
  assign _T_304 = _T_302 | _T_303; // @[Consts.scala 93:41]
  assign _T_305 = s1_req_cmd == 5'h7; // @[Consts.scala 93:65]
  assign _T_306 = _T_304 | _T_305; // @[Consts.scala 93:58]
  assign _T_307 = s1_req_cmd == 5'h4; // @[package.scala 14:47]
  assign _T_308 = s1_req_cmd == 5'h9; // @[package.scala 14:47]
  assign _T_311 = _T_307 | _T_308; // @[package.scala 14:62]
  assign _T_309 = s1_req_cmd == 5'ha; // @[package.scala 14:47]
  assign _T_312 = _T_311 | _T_309; // @[package.scala 14:62]
  assign _T_310 = s1_req_cmd == 5'hb; // @[package.scala 14:47]
  assign _T_313 = _T_312 | _T_310; // @[package.scala 14:62]
  assign _T_314 = s1_req_cmd == 5'h8; // @[package.scala 14:47]
  assign _T_315 = s1_req_cmd == 5'hc; // @[package.scala 14:47]
  assign _T_319 = _T_314 | _T_315; // @[package.scala 14:62]
  assign _T_316 = s1_req_cmd == 5'hd; // @[package.scala 14:47]
  assign _T_320 = _T_319 | _T_316; // @[package.scala 14:62]
  assign _T_317 = s1_req_cmd == 5'he; // @[package.scala 14:47]
  assign _T_321 = _T_320 | _T_317; // @[package.scala 14:62]
  assign _T_318 = s1_req_cmd == 5'hf; // @[package.scala 14:47]
  assign _T_322 = _T_321 | _T_318; // @[package.scala 14:62]
  assign _T_323 = _T_313 | _T_322; // @[Consts.scala 91:44]
  assign s1_read = _T_306 | _T_323; // @[Consts.scala 93:75]
  assign s2_valid_masked = s2_valid & _T_738; // @[DCache.scala 234:34]
  assign _T_749 = s2_req_cmd == 5'h0; // @[Consts.scala 93:31]
  assign _T_750 = s2_req_cmd == 5'h6; // @[Consts.scala 93:48]
  assign _T_751 = _T_749 | _T_750; // @[Consts.scala 93:41]
  assign _T_752 = s2_req_cmd == 5'h7; // @[Consts.scala 93:65]
  assign _T_753 = _T_751 | _T_752; // @[Consts.scala 93:58]
  assign _T_754 = s2_req_cmd == 5'h4; // @[package.scala 14:47]
  assign _T_755 = s2_req_cmd == 5'h9; // @[package.scala 14:47]
  assign _T_758 = _T_754 | _T_755; // @[package.scala 14:62]
  assign _T_756 = s2_req_cmd == 5'ha; // @[package.scala 14:47]
  assign _T_759 = _T_758 | _T_756; // @[package.scala 14:62]
  assign _T_757 = s2_req_cmd == 5'hb; // @[package.scala 14:47]
  assign _T_760 = _T_759 | _T_757; // @[package.scala 14:62]
  assign _T_761 = s2_req_cmd == 5'h8; // @[package.scala 14:47]
  assign _T_762 = s2_req_cmd == 5'hc; // @[package.scala 14:47]
  assign _T_766 = _T_761 | _T_762; // @[package.scala 14:62]
  assign _T_763 = s2_req_cmd == 5'hd; // @[package.scala 14:47]
  assign _T_767 = _T_766 | _T_763; // @[package.scala 14:62]
  assign _T_764 = s2_req_cmd == 5'he; // @[package.scala 14:47]
  assign _T_768 = _T_767 | _T_764; // @[package.scala 14:62]
  assign _T_765 = s2_req_cmd == 5'hf; // @[package.scala 14:47]
  assign _T_769 = _T_768 | _T_765; // @[package.scala 14:62]
  assign _T_770 = _T_760 | _T_769; // @[Consts.scala 91:44]
  assign s2_read = _T_753 | _T_770; // @[Consts.scala 93:75]
  assign _T_771 = s2_req_cmd == 5'h1; // @[Consts.scala 94:32]
  assign _T_772 = s2_req_cmd == 5'h11; // @[Consts.scala 94:49]
  assign _T_773 = _T_771 | _T_772; // @[Consts.scala 94:42]
  assign _T_775 = _T_773 | _T_752; // @[Consts.scala 94:59]
  assign s2_write = _T_775 | _T_770; // @[Consts.scala 94:76]
  assign s2_readwrite = s2_read | s2_write; // @[DCache.scala 247:30]
  assign _T_1033 = s2_valid_masked & s2_readwrite; // @[DCache.scala 282:51]
  assign _T_926 = s2_req_cmd == 5'h3; // @[Consts.scala 95:54]
  assign _T_927 = s2_write | _T_926; // @[Consts.scala 95:47]
  assign _T_929 = _T_927 | _T_750; // @[Consts.scala 95:64]
  assign _T_931 = {s2_write,_T_929,s2_hit_state_state}; // @[Cat.scala 30:58]
  assign _T_989 = 4'h3 == _T_931; // @[Misc.scala 51:20]
  assign _T_986 = 4'h2 == _T_931; // @[Misc.scala 51:20]
  assign _T_983 = 4'h1 == _T_931; // @[Misc.scala 51:20]
  assign _T_980 = 4'h7 == _T_931; // @[Misc.scala 51:20]
  assign _T_977 = 4'h6 == _T_931; // @[Misc.scala 51:20]
  assign _T_974 = 4'hf == _T_931; // @[Misc.scala 51:20]
  assign _T_971 = 4'he == _T_931; // @[Misc.scala 51:20]
  assign _T_968 = 4'h0 == _T_931; // @[Misc.scala 51:20]
  assign _T_965 = 4'h5 == _T_931; // @[Misc.scala 51:20]
  assign _T_962 = 4'h4 == _T_931; // @[Misc.scala 51:20]
  assign _T_959 = 4'hd == _T_931; // @[Misc.scala 51:20]
  assign _T_956 = 4'hc == _T_931; // @[Misc.scala 51:20]
  assign _T_975 = _T_974 | _T_971; // @[Misc.scala 37:9]
  assign _T_978 = _T_977 | _T_975; // @[Misc.scala 37:9]
  assign _T_981 = _T_980 | _T_978; // @[Misc.scala 37:9]
  assign _T_984 = _T_983 | _T_981; // @[Misc.scala 37:9]
  assign _T_987 = _T_986 | _T_984; // @[Misc.scala 37:9]
  assign s2_hit = _T_989 | _T_987; // @[Misc.scala 37:9]
  assign s2_valid_hit_pre_data_ecc = _T_1033 & s2_hit; // @[DCache.scala 282:85]
  assign _T_1417 = s2_valid_hit_pre_data_ecc & s2_write; // @[DCache.scala 345:46]
  assign lrscAddrMatch = lrscAddr == s2_req_addr[39:6]; // @[DCache.scala 331:32]
  assign _T_1255 = lrscValid & lrscAddrMatch; // @[DCache.scala 332:41]
  assign s2_sc_fail = _T_752 & ~_T_1255; // @[DCache.scala 332:26]
  assign _T_1419 = _T_1417 & ~s2_sc_fail; // @[DCache.scala 345:58]
  assign pstore1_valid_pre_kill = _T_1419 | pstore1_held; // @[DCache.scala 361:56]
  assign _T_1591 = pstore1_addr[11:3] == s1_req_addr[11:3]; // @[DCache.scala 414:31]
  assign _T_324 = s1_req_cmd == 5'h1; // @[Consts.scala 94:32]
  assign _T_325 = s1_req_cmd == 5'h11; // @[Consts.scala 94:49]
  assign _T_326 = _T_324 | _T_325; // @[Consts.scala 94:42]
  assign _T_328 = _T_326 | _T_305; // @[Consts.scala 94:59]
  assign s1_write = _T_328 | _T_323; // @[Consts.scala 94:76]
  assign _T_1614 = {pstore1_mask[7],pstore1_mask[6],pstore1_mask[5],pstore1_mask[4],pstore1_mask[3],pstore1_mask[2],pstore1_mask[1],pstore1_mask[0]}; // @[Cat.scala 30:58]
  assign _T_1629 = {_T_1614[7],_T_1614[6],_T_1614[5],_T_1614[4],_T_1614[3],_T_1614[2],_T_1614[1],_T_1614[0]}; // @[Cat.scala 30:58]
  assign _T_701 = s1_req_typ[1:0] >= 2'h1; // @[AMOALU.scala 17:57]
  assign _T_703 = s1_req_addr[0] | _T_701; // @[AMOALU.scala 17:46]
  assign _T_705 = s1_req_addr[0] ? 1'h0 : 1'h1; // @[AMOALU.scala 18:22]
  assign _T_706 = {_T_703,_T_705}; // @[Cat.scala 30:58]
  assign _T_708 = s1_req_addr[1] ? _T_706 : 2'h0; // @[AMOALU.scala 17:22]
  assign _T_709 = s1_req_typ[1:0] >= 2'h2; // @[AMOALU.scala 17:57]
  assign _T_710 = _T_709 ? 2'h3 : 2'h0; // @[AMOALU.scala 17:51]
  assign _T_711 = _T_708 | _T_710; // @[AMOALU.scala 17:46]
  assign _T_713 = s1_req_addr[1] ? 2'h0 : _T_706; // @[AMOALU.scala 18:22]
  assign _T_714 = {_T_711,_T_713}; // @[Cat.scala 30:58]
  assign _T_716 = s1_req_addr[2] ? _T_714 : 4'h0; // @[AMOALU.scala 17:22]
  assign _T_717 = s1_req_typ[1:0] >= 2'h3; // @[AMOALU.scala 17:57]
  assign _T_718 = _T_717 ? 4'hf : 4'h0; // @[AMOALU.scala 17:51]
  assign _T_719 = _T_716 | _T_718; // @[AMOALU.scala 17:46]
  assign _T_721 = s1_req_addr[2] ? 4'h0 : _T_714; // @[AMOALU.scala 18:22]
  assign _T_722 = {_T_719,_T_721}; // @[Cat.scala 30:58]
  assign s1_mask = _T_325 ? 8'h0 : _T_722; // @[DCache.scala 228:20]
  assign _T_1652 = {s1_mask[7],s1_mask[6],s1_mask[5],s1_mask[4],s1_mask[3],s1_mask[2],s1_mask[1],s1_mask[0]}; // @[Cat.scala 30:58]
  assign _T_1667 = {_T_1652[7],_T_1652[6],_T_1652[5],_T_1652[4],_T_1652[3],_T_1652[2],_T_1652[1],_T_1652[0]}; // @[Cat.scala 30:58]
  assign _T_1668 = _T_1629 & _T_1667; // @[DCache.scala 415:38]
  assign _T_1669 = _T_1668 != 8'h0; // @[DCache.scala 415:62]
  assign _T_1670 = pstore1_mask & s1_mask; // @[DCache.scala 415:73]
  assign _T_1671 = _T_1670 != 8'h0; // @[DCache.scala 415:84]
  assign _T_1672 = s1_write ? _T_1669 : _T_1671; // @[DCache.scala 415:8]
  assign _T_1673 = _T_1591 & _T_1672; // @[DCache.scala 414:68]
  assign _T_1674 = pstore1_valid_pre_kill & _T_1673; // @[DCache.scala 417:29]
  assign _T_1677 = pstore2_addr[11:3] == s1_req_addr[11:3]; // @[DCache.scala 414:31]
  assign _T_1700 = {mask[7],mask[6],mask[5],mask[4],mask[3],mask[2],mask[1],mask[0]}; // @[Cat.scala 30:58]
  assign _T_1715 = {_T_1700[7],_T_1700[6],_T_1700[5],_T_1700[4],_T_1700[3],_T_1700[2],_T_1700[1],_T_1700[0]}; // @[Cat.scala 30:58]
  assign _T_1754 = _T_1715 & _T_1667; // @[DCache.scala 415:38]
  assign _T_1755 = _T_1754 != 8'h0; // @[DCache.scala 415:62]
  assign _T_1756 = mask & s1_mask; // @[DCache.scala 415:73]
  assign _T_1757 = _T_1756 != 8'h0; // @[DCache.scala 415:84]
  assign _T_1758 = s1_write ? _T_1755 : _T_1757; // @[DCache.scala 415:8]
  assign _T_1759 = _T_1677 & _T_1758; // @[DCache.scala 414:68]
  assign _T_1760 = pstore2_valid & _T_1759; // @[DCache.scala 418:21]
  assign s1_hazard = _T_1674 | _T_1760; // @[DCache.scala 417:71]
  assign s1_raw_hazard = s1_read & s1_hazard; // @[DCache.scala 419:31]
  assign _T_1761 = s1_valid & s1_raw_hazard; // @[DCache.scala 424:18]
  assign _T_958 = _T_956 ? 2'h1 : 2'h0; // @[Misc.scala 37:36]
  assign _T_961 = _T_959 ? 2'h2 : _T_958; // @[Misc.scala 37:36]
  assign _T_964 = _T_962 ? 2'h1 : _T_961; // @[Misc.scala 37:36]
  assign _T_967 = _T_965 ? 2'h2 : _T_964; // @[Misc.scala 37:36]
  assign _T_970 = _T_968 ? 2'h0 : _T_967; // @[Misc.scala 37:36]
  assign _T_973 = _T_971 ? 2'h3 : _T_970; // @[Misc.scala 37:36]
  assign _T_976 = _T_974 ? 2'h3 : _T_973; // @[Misc.scala 37:36]
  assign _T_979 = _T_977 ? 2'h2 : _T_976; // @[Misc.scala 37:36]
  assign _T_982 = _T_980 ? 2'h3 : _T_979; // @[Misc.scala 37:36]
  assign _T_985 = _T_983 ? 2'h1 : _T_982; // @[Misc.scala 37:36]
  assign _T_988 = _T_986 ? 2'h2 : _T_985; // @[Misc.scala 37:36]
  assign s2_grow_param = _T_989 ? 2'h3 : _T_988; // @[Misc.scala 37:36]
  assign _T_1195 = s2_hit_state_state == s2_grow_param; // @[Metadata.scala 46:46]
  assign s2_update_meta = ~_T_1195; // @[Metadata.scala 47:40]
  assign _T_1201 = s2_valid_hit_pre_data_ecc & s2_update_meta; // @[DCache.scala 301:41]
  assign _T_1202 = io_cpu_s2_nack | _T_1201; // @[DCache.scala 301:24]
  assign s1_readwrite = s1_read | s1_write; // @[DCache.scala 146:30]
  assign _T_543 = s1_valid & s1_readwrite; // @[DCache.scala 193:18]
  assign _T_544 = _T_543 & tlb_io_resp_miss; // @[DCache.scala 193:34]
  assign _GEN_74 = _T_1202 | _T_544; // @[DCache.scala 301:61]
  assign _GEN_98 = _T_1761 | _GEN_74; // @[DCache.scala 424:36]
  assign _GEN_219 = probeNack | _GEN_98; // @[DCache.scala 635:24]
  assign s1_nack = s2_probe ? _GEN_219 : _GEN_98; // @[DCache.scala 620:21]
  assign s1_valid_not_nacked = s1_valid & ~s1_nack; // @[DCache.scala 136:38]
  assign s0_clk_en = metaArb_io_out_valid & ~metaArb_io_out_bits_write; // @[DCache.scala 138:40]
  assign _T_300 = {metaArb_io_out_bits_addr[39:6],io_cpu_req_bits_addr[5:0]}; // @[Cat.scala 30:58]
  assign _GEN_9 = ~metaArb_io_in_7_ready | io_cpu_req_bits_phys; // @[DCache.scala 142:36]
  assign s1_sfence = s1_req_cmd == 5'h14; // @[DCache.scala 147:30]
  assign can_acquire_before_release = ~release_ack_wait; // @[DCache.scala 154:36]
  assign inWriteback = _T_3315 | _T_3314; // @[package.scala 14:62]
  assign _T_357 = release_state == 3'h0; // @[DCache.scala 159:38]
  assign _T_359 = _T_357 & ~cached_grant_wait; // @[DCache.scala 159:51]
  assign _T_361 = _T_359 & ~s1_nack; // @[DCache.scala 159:73]
  assign _T_388 = io_cpu_req_bits_cmd == 5'h0; // @[Consts.scala 93:31]
  assign _T_389 = io_cpu_req_bits_cmd == 5'h6; // @[Consts.scala 93:48]
  assign _T_390 = _T_388 | _T_389; // @[Consts.scala 93:41]
  assign _T_391 = io_cpu_req_bits_cmd == 5'h7; // @[Consts.scala 93:65]
  assign _T_392 = _T_390 | _T_391; // @[Consts.scala 93:58]
  assign _T_393 = io_cpu_req_bits_cmd == 5'h4; // @[package.scala 14:47]
  assign _T_394 = io_cpu_req_bits_cmd == 5'h9; // @[package.scala 14:47]
  assign _T_395 = io_cpu_req_bits_cmd == 5'ha; // @[package.scala 14:47]
  assign _T_396 = io_cpu_req_bits_cmd == 5'hb; // @[package.scala 14:47]
  assign _T_397 = _T_393 | _T_394; // @[package.scala 14:62]
  assign _T_398 = _T_397 | _T_395; // @[package.scala 14:62]
  assign _T_399 = _T_398 | _T_396; // @[package.scala 14:62]
  assign _T_400 = io_cpu_req_bits_cmd == 5'h8; // @[package.scala 14:47]
  assign _T_401 = io_cpu_req_bits_cmd == 5'hc; // @[package.scala 14:47]
  assign _T_402 = io_cpu_req_bits_cmd == 5'hd; // @[package.scala 14:47]
  assign _T_403 = io_cpu_req_bits_cmd == 5'he; // @[package.scala 14:47]
  assign _T_404 = io_cpu_req_bits_cmd == 5'hf; // @[package.scala 14:47]
  assign _T_405 = _T_400 | _T_401; // @[package.scala 14:62]
  assign _T_406 = _T_405 | _T_402; // @[package.scala 14:62]
  assign _T_407 = _T_406 | _T_403; // @[package.scala 14:62]
  assign _T_408 = _T_407 | _T_404; // @[package.scala 14:62]
  assign _T_409 = _T_399 | _T_408; // @[Consts.scala 91:44]
  assign s0_read = _T_392 | _T_409; // @[Consts.scala 93:75]
  assign _T_410 = io_cpu_req_bits_cmd == 5'h1; // @[package.scala 14:47]
  assign _T_411 = io_cpu_req_bits_cmd == 5'h3; // @[package.scala 14:47]
  assign _T_412 = _T_410 | _T_411; // @[package.scala 14:62]
  assign res = ~_T_412; // @[DCache.scala 912:15]
  assign _T_440 = io_cpu_req_bits_cmd == 5'h11; // @[Consts.scala 94:49]
  assign _T_441 = _T_410 | _T_440; // @[Consts.scala 94:42]
  assign _T_443 = _T_441 | _T_391; // @[Consts.scala 94:59]
  assign _T_461 = _T_443 | _T_409; // @[Consts.scala 94:76]
  assign _T_466 = _T_461 & _T_440; // @[DCache.scala 918:23]
  assign _T_467 = s0_read | _T_466; // @[DCache.scala 917:21]
  assign _T_469 = ~_T_467 | res; // @[DCache.scala 913:28]
  assign _T_471 = _T_469 | reset; // @[DCache.scala 913:11]
  assign _T_473 = io_cpu_req_valid & res; // @[DCache.scala 167:46]
  assign _T_477 = ~dataArb_io_in_3_ready & s0_read; // @[DCache.scala 173:33]
  assign _GEN_16 = _T_477 ? 1'h0 : _T_361; // @[DCache.scala 173:45]
  assign _GEN_18 = metaArb_io_in_7_ready ? _GEN_16 : 1'h0; // @[DCache.scala 181:34]
  assign _T_540 = ~tlb_io_req_ready & ~tlb_io_ptw_resp_valid; // @[DCache.scala 192:27]
  assign _T_542 = _T_540 & ~io_cpu_req_bits_phys; // @[DCache.scala 192:53]
  assign _GEN_19 = _T_542 ? 1'h0 : _GEN_18; // @[DCache.scala 192:79]
  assign s1_victim_way = lfsr[1:0]; // @[Replacement.scala 19:44]
  assign _T_600 = tag_array_0_s1_meta_data;
  assign _T_607 = tag_array_1_s1_meta_data;
  assign _T_614 = tag_array_2_s1_meta_data;
  assign _T_621 = tag_array_3_s1_meta_data;
  assign s1_tag = tlb_io_resp_paddr[31:12]; // @[DCache.scala 219:29]
  assign _T_624 = _T_600[21:20] > 2'h0; // @[Metadata.scala 50:45]
  assign _T_625 = _T_600[19:0] == s1_tag; // @[DCache.scala 220:83]
  assign _T_626 = _T_624 & _T_625; // @[DCache.scala 220:74]
  assign _T_627 = _T_607[21:20] > 2'h0; // @[Metadata.scala 50:45]
  assign _T_628 = _T_607[19:0] == s1_tag; // @[DCache.scala 220:83]
  assign _T_629 = _T_627 & _T_628; // @[DCache.scala 220:74]
  assign _T_630 = _T_614[21:20] > 2'h0; // @[Metadata.scala 50:45]
  assign _T_631 = _T_614[19:0] == s1_tag; // @[DCache.scala 220:83]
  assign _T_632 = _T_630 & _T_631; // @[DCache.scala 220:74]
  assign _T_633 = _T_621[21:20] > 2'h0; // @[Metadata.scala 50:45]
  assign _T_634 = _T_621[19:0] == s1_tag; // @[DCache.scala 220:83]
  assign _T_635 = _T_633 & _T_634; // @[DCache.scala 220:74]
  assign s1_meta_hit_way = {_T_635,_T_632,_T_629,_T_626}; // @[Cat.scala 30:58]
  assign _T_642 = _T_625 & ~s1_flush_valid; // @[DCache.scala 222:59]
  assign _T_643 = _T_642 ? _T_600[21:20] : 2'h0; // @[DCache.scala 222:41]
  assign _T_646 = _T_628 & ~s1_flush_valid; // @[DCache.scala 222:59]
  assign _T_647 = _T_646 ? _T_607[21:20] : 2'h0; // @[DCache.scala 222:41]
  assign _T_650 = _T_631 & ~s1_flush_valid; // @[DCache.scala 222:59]
  assign _T_651 = _T_650 ? _T_614[21:20] : 2'h0; // @[DCache.scala 222:41]
  assign _T_654 = _T_634 & ~s1_flush_valid; // @[DCache.scala 222:59]
  assign _T_655 = _T_654 ? _T_621[21:20] : 2'h0; // @[DCache.scala 222:41]
  assign _T_656 = _T_643 | _T_647; // @[DCache.scala 223:19]
  assign _T_657 = _T_656 | _T_651; // @[DCache.scala 223:19]
  assign s1_meta_hit_state_state = _T_657 | _T_655; // @[DCache.scala 223:19]
  assign _T_665 = s1_victim_way == 2'h1; // @[package.scala 31:81]
  assign _T_667 = s1_victim_way == 2'h2; // @[package.scala 31:81]
  assign _T_669 = s1_victim_way == 2'h3; // @[package.scala 31:81]
  assign s2_hit_valid = s2_hit_state_state > 2'h0; // @[Metadata.scala 50:45]
  assign _T_1061 = 4'h1 << _T_1060; // @[OneHot.scala 45:35]
  assign s2_victim_way = s2_hit_valid ? s2_hit_way : _T_1061; // @[DCache.scala 292:26]
  assign releaseWay = _T_3317 ? s2_victim_way : s2_probe_way; // @[DCache.scala 659:81]
  assign _T_670 = inWriteback ? releaseWay : s1_meta_hit_way; // @[DCache.scala 226:61]
  assign s1_all_data_ways_4 = {auto_out_d_bits_data[63:56],auto_out_d_bits_data[55:48],auto_out_d_bits_data[47:40],auto_out_d_bits_data[39:32],auto_out_d_bits_data[31:24],auto_out_d_bits_data[23:16],auto_out_d_bits_data[15:8],auto_out_d_bits_data[7:0]}; // @[Cat.scala 30:58]
  assign _T_724 = s1_valid_masked & ~s1_sfence; // @[DCache.scala 230:52]
  assign _T_742 = s1_valid_not_nacked | s1_flush_valid; // @[DCache.scala 239:29]
  assign s2_vaddr = {_T_746[39:12],s2_req_addr[11:0]}; // @[Cat.scala 30:58]
  assign en = s1_valid | inWriteback; // @[DCache.scala 258:23]
  assign _T_3079 = auto_out_d_bits_opcode == 3'h0; // @[package.scala 14:47]
  assign _T_3081 = grantIsUncachedData | _T_3079; // @[package.scala 14:62]
  assign _T_3080 = auto_out_d_bits_opcode == 3'h2; // @[package.scala 14:47]
  assign grantIsUncached = _T_3081 | _T_3080; // @[package.scala 14:62]
  assign _GEN_129 = grantIsUncachedData ? 5'h10 : {{1'd0}, _T_670}; // @[DCache.scala 516:34]
  assign _GEN_137 = grantIsUncached ? _GEN_129 : {{1'd0}, _T_670}; // @[DCache.scala 507:35]
  assign _GEN_149 = grantIsCached ? {{1'd0}, _T_670} : _GEN_137; // @[DCache.scala 498:26]
  assign s1_data_way = _T_3094 ? _GEN_149 : {{1'd0}, _T_670}; // @[DCache.scala 497:26]
  assign s1_all_data_ways_0 = data_io_resp_0; // @[DCache.scala 227:29 DCache.scala 227:29]
  assign _T_859 = s1_data_way[0] ? s1_all_data_ways_0 : 64'h0; // @[Mux.scala 19:72]
  assign s1_all_data_ways_1 = data_io_resp_1; // @[DCache.scala 227:29 DCache.scala 227:29]
  assign _T_860 = s1_data_way[1] ? s1_all_data_ways_1 : 64'h0; // @[Mux.scala 19:72]
  assign s1_all_data_ways_2 = data_io_resp_2; // @[DCache.scala 227:29 DCache.scala 227:29]
  assign _T_861 = s1_data_way[2] ? s1_all_data_ways_2 : 64'h0; // @[Mux.scala 19:72]
  assign s1_all_data_ways_3 = data_io_resp_3; // @[DCache.scala 227:29 DCache.scala 227:29]
  assign _T_862 = s1_data_way[3] ? s1_all_data_ways_3 : 64'h0; // @[Mux.scala 19:72]
  assign _T_863 = s1_data_way[4] ? s1_all_data_ways_4 : 64'h0; // @[Mux.scala 19:72]
  assign _T_864 = _T_859 | _T_860; // @[Mux.scala 19:72]
  assign _T_865 = _T_864 | _T_861; // @[Mux.scala 19:72]
  assign _T_866 = _T_865 | _T_862; // @[Mux.scala 19:72]
  assign _T_867 = _T_866 | _T_863; // @[Mux.scala 19:72]
  assign _T_871 = en | _T_3094; // @[DCache.scala 264:58]
  assign _T_1023 = {s2_data[31:24],s2_data[23:16],s2_data[15:8],s2_data[7:0]}; // @[Cat.scala 30:58]
  assign _T_1026 = {s2_data[63:56],s2_data[55:48],s2_data[47:40],s2_data[39:32]}; // @[Cat.scala 30:58]
  assign s2_data_corrected = {s2_data[63:56],s2_data[55:48],s2_data[47:40],s2_data[39:32],s2_data[31:24],s2_data[23:16],s2_data[15:8],s2_data[7:0]}; // @[Cat.scala 30:58]
  assign _T_1045 = _T_1033 & ~s2_hit; // @[DCache.scala 285:73]
  assign s2_valid_miss = _T_1045 & can_acquire_before_release; // @[DCache.scala 285:84]
  assign _T_1047 = s2_valid_miss & ~s2_uncached; // @[DCache.scala 286:44]
  assign s2_valid_cached_miss = _T_1047 & ~uncachedInFlight_0; // @[DCache.scala 286:60]
  assign s2_want_victimize = s2_valid_cached_miss | s2_flush_valid_pre_tag_ecc; // @[DCache.scala 288:102]
  assign _T_1054 = s2_valid_miss & s2_uncached; // @[DCache.scala 291:49]
  assign s2_valid_uncached_pending = _T_1054 & ~uncachedInFlight_0; // @[DCache.scala 291:64]
  assign s2_victim_state_state = s2_hit_valid ? s2_hit_state_state : _T_1068_state; // @[DCache.scala 294:28]
  assign _T_1084 = _T_1082 ? 3'h5 : 3'h0; // @[Misc.scala 40:36]
  assign _T_1088 = _T_1086 ? 3'h2 : _T_1084; // @[Misc.scala 40:36]
  assign _T_1092 = _T_1090 ? 3'h1 : _T_1088; // @[Misc.scala 40:36]
  assign _T_1096 = _T_1094 ? 3'h1 : _T_1092; // @[Misc.scala 40:36]
  assign _T_1100 = _T_1098 ? 3'h2 : _T_1096; // @[Misc.scala 40:36]
  assign _T_1104 = _T_1102 ? 3'h4 : _T_1100; // @[Misc.scala 40:36]
  assign _T_1105 = _T_1102 ? 2'h1 : 2'h0; // @[Misc.scala 40:63]
  assign _T_1108 = _T_1106 ? 3'h0 : _T_1104; // @[Misc.scala 40:36]
  assign _T_1109 = _T_1106 ? 2'h1 : _T_1105; // @[Misc.scala 40:63]
  assign _T_1112 = _T_1110 ? 3'h0 : _T_1108; // @[Misc.scala 40:36]
  assign _T_1113 = _T_1110 ? 2'h1 : _T_1109; // @[Misc.scala 40:63]
  assign _T_1116 = _T_1114 ? 3'h5 : _T_1112; // @[Misc.scala 40:36]
  assign _T_1117 = _T_1114 ? 2'h0 : _T_1113; // @[Misc.scala 40:63]
  assign _T_1120 = _T_1118 ? 3'h4 : _T_1116; // @[Misc.scala 40:36]
  assign _T_1121 = _T_1118 ? 2'h1 : _T_1117; // @[Misc.scala 40:63]
  assign _T_1124 = _T_1122 ? 3'h3 : _T_1120; // @[Misc.scala 40:36]
  assign _T_1125 = _T_1122 ? 2'h2 : _T_1121; // @[Misc.scala 40:63]
  assign s2_report_param = _T_1126 ? 3'h3 : _T_1124; // @[Misc.scala 40:36]
  assign probeNewCoh_state = _T_1126 ? 2'h2 : _T_1125; // @[Misc.scala 40:63]
  assign _T_1135 = {2'h2,s2_victim_state_state}; // @[Cat.scala 30:58]
  assign _T_1148 = 4'h8 == _T_1135; // @[Misc.scala 58:20]
  assign _T_1150 = _T_1148 ? 3'h5 : 3'h0; // @[Misc.scala 40:36]
  assign _T_1152 = 4'h9 == _T_1135; // @[Misc.scala 58:20]
  assign _T_1154 = _T_1152 ? 3'h2 : _T_1150; // @[Misc.scala 40:36]
  assign _T_1156 = 4'ha == _T_1135; // @[Misc.scala 58:20]
  assign _T_1158 = _T_1156 ? 3'h1 : _T_1154; // @[Misc.scala 40:36]
  assign _T_1160 = 4'hb == _T_1135; // @[Misc.scala 58:20]
  assign _T_1162 = _T_1160 ? 3'h1 : _T_1158; // @[Misc.scala 40:36]
  assign _T_1164 = 4'h4 == _T_1135; // @[Misc.scala 58:20]
  assign _T_1165 = _T_1164 ? 1'h0 : _T_1160; // @[Misc.scala 40:9]
  assign _T_1166 = _T_1164 ? 3'h2 : _T_1162; // @[Misc.scala 40:36]
  assign _T_1168 = 4'h5 == _T_1135; // @[Misc.scala 58:20]
  assign _T_1169 = _T_1168 ? 1'h0 : _T_1165; // @[Misc.scala 40:9]
  assign _T_1170 = _T_1168 ? 3'h4 : _T_1166; // @[Misc.scala 40:36]
  assign _T_1171 = _T_1168 ? 2'h1 : 2'h0; // @[Misc.scala 40:63]
  assign _T_1172 = 4'h6 == _T_1135; // @[Misc.scala 58:20]
  assign _T_1173 = _T_1172 ? 1'h0 : _T_1169; // @[Misc.scala 40:9]
  assign _T_1174 = _T_1172 ? 3'h0 : _T_1170; // @[Misc.scala 40:36]
  assign _T_1175 = _T_1172 ? 2'h1 : _T_1171; // @[Misc.scala 40:63]
  assign _T_1176 = 4'h7 == _T_1135; // @[Misc.scala 58:20]
  assign _T_1177 = _T_1176 | _T_1173; // @[Misc.scala 40:9]
  assign _T_1178 = _T_1176 ? 3'h0 : _T_1174; // @[Misc.scala 40:36]
  assign _T_1179 = _T_1176 ? 2'h1 : _T_1175; // @[Misc.scala 40:63]
  assign _T_1180 = 4'h0 == _T_1135; // @[Misc.scala 58:20]
  assign _T_1181 = _T_1180 ? 1'h0 : _T_1177; // @[Misc.scala 40:9]
  assign _T_1182 = _T_1180 ? 3'h5 : _T_1178; // @[Misc.scala 40:36]
  assign _T_1183 = _T_1180 ? 2'h0 : _T_1179; // @[Misc.scala 40:63]
  assign _T_1184 = 4'h1 == _T_1135; // @[Misc.scala 58:20]
  assign _T_1185 = _T_1184 ? 1'h0 : _T_1181; // @[Misc.scala 40:9]
  assign _T_1186 = _T_1184 ? 3'h4 : _T_1182; // @[Misc.scala 40:36]
  assign _T_1187 = _T_1184 ? 2'h1 : _T_1183; // @[Misc.scala 40:63]
  assign _T_1188 = 4'h2 == _T_1135; // @[Misc.scala 58:20]
  assign _T_1189 = _T_1188 ? 1'h0 : _T_1185; // @[Misc.scala 40:9]
  assign _T_1190 = _T_1188 ? 3'h3 : _T_1186; // @[Misc.scala 40:36]
  assign _T_1191 = _T_1188 ? 2'h2 : _T_1187; // @[Misc.scala 40:63]
  assign _T_1192 = 4'h3 == _T_1135; // @[Misc.scala 58:20]
  assign s2_victim_dirty = _T_1192 | _T_1189; // @[Misc.scala 40:9]
  assign s2_shrink_param = _T_1192 ? 3'h3 : _T_1190; // @[Misc.scala 40:36]
  assign voluntaryNewCoh_state = _T_1192 ? 2'h2 : _T_1191; // @[Misc.scala 40:63]
  assign _T_1197 = s2_valid & ~s2_valid_hit_pre_data_ecc; // @[DCache.scala 300:30]
  assign _T_1198 = s2_valid_uncached_pending & auto_out_a_ready; // @[DCache.scala 300:78]
  assign _T_1200 = _T_1197 & ~_T_1198; // @[DCache.scala 300:47]
  assign _T_1234 = s2_want_victimize & ~s2_victim_dirty; // @[DCache.scala 317:84]
  assign _T_1244_state = s2_valid_hit_pre_data_ecc ? s2_grow_param : 2'h0; // @[DCache.scala 322:82]
  assign _T_1251 = lrscCount > 7'h0; // @[DCache.scala 329:34]
  assign lrscBackingOff = _T_1251 & ~lrscValid; // @[DCache.scala 329:38]
  assign _T_1257 = s2_valid_hit_pre_data_ecc & _T_750; // @[DCache.scala 333:23]
  assign _T_1259 = _T_1257 & ~cached_grant_wait; // @[DCache.scala 333:32]
  assign _T_1260 = _T_1259 | s2_valid_cached_miss; // @[DCache.scala 333:54]
  assign _T_1268 = lrscCount - 7'h1; // @[DCache.scala 337:49]
  assign _T_1269 = s2_valid_masked & lrscValid; // @[DCache.scala 338:29]
  assign _T_1278 = s1_valid_not_nacked & s1_write; // @[DCache.scala 347:63]
  assign _T_1339 = s1_write & _T_325; // @[DCache.scala 918:23]
  assign _T_1340 = s1_read | _T_1339; // @[DCache.scala 917:21]
  assign _T_1344 = s2_valid & s2_write; // @[DCache.scala 354:39]
  assign pstore_drain_opportunistic = ~_T_473; // @[DCache.scala 357:36]
  assign pstore1_valid_likely = _T_1344 | pstore1_held; // @[DCache.scala 360:51]
  assign _T_1426 = pstore1_valid_likely & pstore2_valid; // @[DCache.scala 365:54]
  assign _T_1427 = s1_valid & s1_write; // @[DCache.scala 365:85]
  assign _T_1428 = _T_1427 | pstore1_rmw; // @[DCache.scala 365:98]
  assign pstore_drain_structural = _T_1426 & _T_1428; // @[DCache.scala 365:71]
  assign _T_1438 = pstore1_valid_pre_kill == pstore1_valid_pre_kill; // @[DCache.scala 366:63]
  assign _T_1439 = pstore1_rmw | _T_1438; // @[DCache.scala 366:22]
  assign _T_1441 = _T_1439 | reset; // @[DCache.scala 366:9]
  assign _T_1457 = pstore1_valid_pre_kill & ~pstore1_rmw; // @[DCache.scala 374:41]
  assign _T_1458 = _T_1457 | pstore2_valid; // @[DCache.scala 374:58]
  assign _T_1459 = pstore_drain_opportunistic | releaseInFlight; // @[DCache.scala 374:107]
  assign _T_1460 = _T_1458 & _T_1459; // @[DCache.scala 374:76]
  assign pstore_drain = pstore_drain_structural | _T_1460; // @[DCache.scala 373:48]
  assign _T_1470 = pstore1_valid_pre_kill & pstore2_valid; // @[DCache.scala 377:71]
  assign _T_1474 = pstore2_valid == pstore_drain; // @[DCache.scala 378:79]
  assign advance_pstore1 = pstore1_valid_pre_kill & _T_1474; // @[DCache.scala 378:61]
  assign _T_1476 = pstore2_valid & ~pstore_drain; // @[DCache.scala 379:34]
  assign pstore1_storegen_data = amoalu_io_out; // @[DCache.scala 748:27]
  assign pstore2_storegen_data = {_T_1529,_T_1523,_T_1517,_T_1511,_T_1505,_T_1499,_T_1493,_T_1487}; // @[Cat.scala 30:58]
  assign _T_1560 = pstore2_valid ? pstore2_addr : pstore1_addr; // @[DCache.scala 405:36]
  assign _T_1565 = pstore2_valid ? mask : pstore1_mask; // @[DCache.scala 410:47]
  assign _T_1584 = {_T_1565[3],_T_1565[2],_T_1565[1],_T_1565[0]}; // @[Cat.scala 30:58]
  assign _T_1587 = {_T_1565[7],_T_1565[6],_T_1565[5],_T_1565[4]}; // @[Cat.scala 30:58]
  assign _T_1765 = {~uncachedInFlight_0, 1'h0}; // @[DCache.scala 430:59]
  assign a_source = _T_1765[0] ? 1'h0 : 1'h1; // @[Mux.scala 31:69]
  assign acquire_address = {s2_req_addr[39:6], 6'h0}; // @[DCache.scala 431:49]
  assign a_size = s2_req_typ[1:0]; // @[Consts.scala 19:28]
  assign _T_1822 = {{1'd0}, a_size}; // @[Misc.scala 206:34]
  assign _T_1824 = 4'h1 << _T_1822[1:0]; // @[OneHot.scala 52:12]
  assign _T_1826 = _T_1824[2:0] | 3'h1; // @[Misc.scala 206:81]
  assign _T_1827 = a_size >= 2'h3; // @[Misc.scala 210:21]
  assign _T_1832 = _T_1826[2] & ~s2_req_addr[2]; // @[Misc.scala 219:38]
  assign _T_1833 = _T_1827 | _T_1832; // @[Misc.scala 219:29]
  assign _T_1835 = _T_1826[2] & s2_req_addr[2]; // @[Misc.scala 219:38]
  assign _T_1836 = _T_1827 | _T_1835; // @[Misc.scala 219:29]
  assign _T_1840 = ~s2_req_addr[2] & ~s2_req_addr[1]; // @[Misc.scala 218:27]
  assign _T_1841 = _T_1826[1] & _T_1840; // @[Misc.scala 219:38]
  assign _T_1842 = _T_1833 | _T_1841; // @[Misc.scala 219:29]
  assign _T_1843 = ~s2_req_addr[2] & s2_req_addr[1]; // @[Misc.scala 218:27]
  assign _T_1844 = _T_1826[1] & _T_1843; // @[Misc.scala 219:38]
  assign _T_1845 = _T_1833 | _T_1844; // @[Misc.scala 219:29]
  assign _T_1846 = s2_req_addr[2] & ~s2_req_addr[1]; // @[Misc.scala 218:27]
  assign _T_1847 = _T_1826[1] & _T_1846; // @[Misc.scala 219:38]
  assign _T_1848 = _T_1836 | _T_1847; // @[Misc.scala 219:29]
  assign _T_1849 = s2_req_addr[2] & s2_req_addr[1]; // @[Misc.scala 218:27]
  assign _T_1850 = _T_1826[1] & _T_1849; // @[Misc.scala 219:38]
  assign _T_1851 = _T_1836 | _T_1850; // @[Misc.scala 219:29]
  assign _T_1855 = _T_1840 & ~s2_req_addr[0]; // @[Misc.scala 218:27]
  assign _T_1856 = _T_1826[0] & _T_1855; // @[Misc.scala 219:38]
  assign _T_1857 = _T_1842 | _T_1856; // @[Misc.scala 219:29]
  assign _T_1858 = _T_1840 & s2_req_addr[0]; // @[Misc.scala 218:27]
  assign _T_1859 = _T_1826[0] & _T_1858; // @[Misc.scala 219:38]
  assign _T_1860 = _T_1842 | _T_1859; // @[Misc.scala 219:29]
  assign _T_1861 = _T_1843 & ~s2_req_addr[0]; // @[Misc.scala 218:27]
  assign _T_1862 = _T_1826[0] & _T_1861; // @[Misc.scala 219:38]
  assign _T_1863 = _T_1845 | _T_1862; // @[Misc.scala 219:29]
  assign _T_1864 = _T_1843 & s2_req_addr[0]; // @[Misc.scala 218:27]
  assign _T_1865 = _T_1826[0] & _T_1864; // @[Misc.scala 219:38]
  assign _T_1866 = _T_1845 | _T_1865; // @[Misc.scala 219:29]
  assign _T_1867 = _T_1846 & ~s2_req_addr[0]; // @[Misc.scala 218:27]
  assign _T_1868 = _T_1826[0] & _T_1867; // @[Misc.scala 219:38]
  assign _T_1869 = _T_1848 | _T_1868; // @[Misc.scala 219:29]
  assign _T_1870 = _T_1846 & s2_req_addr[0]; // @[Misc.scala 218:27]
  assign _T_1871 = _T_1826[0] & _T_1870; // @[Misc.scala 219:38]
  assign _T_1872 = _T_1848 | _T_1871; // @[Misc.scala 219:29]
  assign _T_1873 = _T_1849 & ~s2_req_addr[0]; // @[Misc.scala 218:27]
  assign _T_1874 = _T_1826[0] & _T_1873; // @[Misc.scala 219:38]
  assign _T_1875 = _T_1851 | _T_1874; // @[Misc.scala 219:29]
  assign _T_1876 = _T_1849 & s2_req_addr[0]; // @[Misc.scala 218:27]
  assign _T_1877 = _T_1826[0] & _T_1876; // @[Misc.scala 219:38]
  assign _T_1878 = _T_1851 | _T_1877; // @[Misc.scala 219:29]
  assign get_mask = {_T_1878,_T_1875,_T_1872,_T_1869,_T_1866,_T_1863,_T_1860,_T_1857}; // @[Cat.scala 30:58]
  assign _T_2939 = 5'hf == s2_req_cmd; // @[Mux.scala 46:19]
  assign _T_2940_opcode = _T_2939 ? 3'h2 : 3'h0; // @[Mux.scala 46:16]
  assign _T_2940_param = _T_2939 ? 3'h3 : 3'h0; // @[Mux.scala 46:16]
  assign _T_2874_size = {{2'd0}, a_size}; // @[Edges.scala 476:17 Edges.scala 479:15]
  assign _T_2940_size = _T_2939 ? _T_2874_size : 4'h0; // @[Mux.scala 46:16]
  assign _T_2940_source = _T_2939 & a_source; // @[Mux.scala 46:16]
  assign _T_2940_address = _T_2939 ? s2_req_addr[31:0] : 32'h0; // @[Mux.scala 46:16]
  assign _T_2940_mask = _T_2939 ? get_mask : 8'h0; // @[Mux.scala 46:16]
  assign _T_2940_data = _T_2939 ? pstore1_data : 64'h0; // @[Mux.scala 46:16]
  assign _T_2941 = 5'he == s2_req_cmd; // @[Mux.scala 46:19]
  assign _T_2942_opcode = _T_2941 ? 3'h2 : _T_2940_opcode; // @[Mux.scala 46:16]
  assign _T_2942_param = _T_2941 ? 3'h2 : _T_2940_param; // @[Mux.scala 46:16]
  assign _T_2942_size = _T_2941 ? _T_2874_size : _T_2940_size; // @[Mux.scala 46:16]
  assign _T_2942_source = _T_2941 ? a_source : _T_2940_source; // @[Mux.scala 46:16]
  assign _T_2942_address = _T_2941 ? s2_req_addr[31:0] : _T_2940_address; // @[Mux.scala 46:16]
  assign _T_2942_mask = _T_2941 ? get_mask : _T_2940_mask; // @[Mux.scala 46:16]
  assign _T_2942_data = _T_2941 ? pstore1_data : _T_2940_data; // @[Mux.scala 46:16]
  assign _T_2943 = 5'hd == s2_req_cmd; // @[Mux.scala 46:19]
  assign _T_2944_opcode = _T_2943 ? 3'h2 : _T_2942_opcode; // @[Mux.scala 46:16]
  assign _T_2944_param = _T_2943 ? 3'h1 : _T_2942_param; // @[Mux.scala 46:16]
  assign _T_2944_size = _T_2943 ? _T_2874_size : _T_2942_size; // @[Mux.scala 46:16]
  assign _T_2944_source = _T_2943 ? a_source : _T_2942_source; // @[Mux.scala 46:16]
  assign _T_2944_address = _T_2943 ? s2_req_addr[31:0] : _T_2942_address; // @[Mux.scala 46:16]
  assign _T_2944_mask = _T_2943 ? get_mask : _T_2942_mask; // @[Mux.scala 46:16]
  assign _T_2944_data = _T_2943 ? pstore1_data : _T_2942_data; // @[Mux.scala 46:16]
  assign _T_2945 = 5'hc == s2_req_cmd; // @[Mux.scala 46:19]
  assign _T_2946_opcode = _T_2945 ? 3'h2 : _T_2944_opcode; // @[Mux.scala 46:16]
  assign _T_2946_param = _T_2945 ? 3'h0 : _T_2944_param; // @[Mux.scala 46:16]
  assign _T_2946_size = _T_2945 ? _T_2874_size : _T_2944_size; // @[Mux.scala 46:16]
  assign _T_2946_source = _T_2945 ? a_source : _T_2944_source; // @[Mux.scala 46:16]
  assign _T_2946_address = _T_2945 ? s2_req_addr[31:0] : _T_2944_address; // @[Mux.scala 46:16]
  assign _T_2946_mask = _T_2945 ? get_mask : _T_2944_mask; // @[Mux.scala 46:16]
  assign _T_2946_data = _T_2945 ? pstore1_data : _T_2944_data; // @[Mux.scala 46:16]
  assign _T_2947 = 5'h8 == s2_req_cmd; // @[Mux.scala 46:19]
  assign _T_2948_opcode = _T_2947 ? 3'h2 : _T_2946_opcode; // @[Mux.scala 46:16]
  assign _T_2948_param = _T_2947 ? 3'h4 : _T_2946_param; // @[Mux.scala 46:16]
  assign _T_2948_size = _T_2947 ? _T_2874_size : _T_2946_size; // @[Mux.scala 46:16]
  assign _T_2948_source = _T_2947 ? a_source : _T_2946_source; // @[Mux.scala 46:16]
  assign _T_2948_address = _T_2947 ? s2_req_addr[31:0] : _T_2946_address; // @[Mux.scala 46:16]
  assign _T_2948_mask = _T_2947 ? get_mask : _T_2946_mask; // @[Mux.scala 46:16]
  assign _T_2948_data = _T_2947 ? pstore1_data : _T_2946_data; // @[Mux.scala 46:16]
  assign _T_2949 = 5'hb == s2_req_cmd; // @[Mux.scala 46:19]
  assign _T_2950_opcode = _T_2949 ? 3'h3 : _T_2948_opcode; // @[Mux.scala 46:16]
  assign _T_2950_param = _T_2949 ? 3'h2 : _T_2948_param; // @[Mux.scala 46:16]
  assign _T_2950_size = _T_2949 ? _T_2874_size : _T_2948_size; // @[Mux.scala 46:16]
  assign _T_2950_source = _T_2949 ? a_source : _T_2948_source; // @[Mux.scala 46:16]
  assign _T_2950_address = _T_2949 ? s2_req_addr[31:0] : _T_2948_address; // @[Mux.scala 46:16]
  assign _T_2950_mask = _T_2949 ? get_mask : _T_2948_mask; // @[Mux.scala 46:16]
  assign _T_2950_data = _T_2949 ? pstore1_data : _T_2948_data; // @[Mux.scala 46:16]
  assign _T_2951 = 5'ha == s2_req_cmd; // @[Mux.scala 46:19]
  assign _T_2952_opcode = _T_2951 ? 3'h3 : _T_2950_opcode; // @[Mux.scala 46:16]
  assign _T_2952_param = _T_2951 ? 3'h1 : _T_2950_param; // @[Mux.scala 46:16]
  assign _T_2952_size = _T_2951 ? _T_2874_size : _T_2950_size; // @[Mux.scala 46:16]
  assign _T_2952_source = _T_2951 ? a_source : _T_2950_source; // @[Mux.scala 46:16]
  assign _T_2952_address = _T_2951 ? s2_req_addr[31:0] : _T_2950_address; // @[Mux.scala 46:16]
  assign _T_2952_mask = _T_2951 ? get_mask : _T_2950_mask; // @[Mux.scala 46:16]
  assign _T_2952_data = _T_2951 ? pstore1_data : _T_2950_data; // @[Mux.scala 46:16]
  assign _T_2953 = 5'h9 == s2_req_cmd; // @[Mux.scala 46:19]
  assign _T_2954_opcode = _T_2953 ? 3'h3 : _T_2952_opcode; // @[Mux.scala 46:16]
  assign _T_2954_param = _T_2953 ? 3'h0 : _T_2952_param; // @[Mux.scala 46:16]
  assign _T_2954_size = _T_2953 ? _T_2874_size : _T_2952_size; // @[Mux.scala 46:16]
  assign _T_2954_source = _T_2953 ? a_source : _T_2952_source; // @[Mux.scala 46:16]
  assign _T_2954_address = _T_2953 ? s2_req_addr[31:0] : _T_2952_address; // @[Mux.scala 46:16]
  assign _T_2954_mask = _T_2953 ? get_mask : _T_2952_mask; // @[Mux.scala 46:16]
  assign _T_2954_data = _T_2953 ? pstore1_data : _T_2952_data; // @[Mux.scala 46:16]
  assign _T_2955 = 5'h4 == s2_req_cmd; // @[Mux.scala 46:19]
  assign atomics_opcode = _T_2955 ? 3'h3 : _T_2954_opcode; // @[Mux.scala 46:16]
  assign atomics_param = _T_2955 ? 3'h3 : _T_2954_param; // @[Mux.scala 46:16]
  assign atomics_size = _T_2955 ? _T_2874_size : _T_2954_size; // @[Mux.scala 46:16]
  assign atomics_source = _T_2955 ? a_source : _T_2954_source; // @[Mux.scala 46:16]
  assign atomics_address = _T_2955 ? s2_req_addr[31:0] : _T_2954_address; // @[Mux.scala 46:16]
  assign atomics_mask = _T_2955 ? get_mask : _T_2954_mask; // @[Mux.scala 46:16]
  assign atomics_data = _T_2955 ? pstore1_data : _T_2954_data; // @[Mux.scala 46:16]
  assign _T_2959 = s2_valid_cached_miss & ~s2_victim_dirty; // @[DCache.scala 454:63]
  assign tl_out_a_valid = _T_2959 | s2_valid_uncached_pending; // @[DCache.scala 454:128]
  assign _T_3052_opcode = s2_read ? atomics_opcode : 3'h0; // @[DCache.scala 455:108]
  assign _T_3052_param = s2_read ? atomics_param : 3'h0; // @[DCache.scala 455:108]
  assign _T_3052_size = s2_read ? atomics_size : _T_2874_size; // @[DCache.scala 455:108]
  assign _T_3052_source = s2_read ? atomics_source : a_source; // @[DCache.scala 455:108]
  assign _T_3052_address = s2_read ? atomics_address : s2_req_addr[31:0]; // @[DCache.scala 455:108]
  assign _T_3052_mask = s2_read ? atomics_mask : get_mask; // @[DCache.scala 455:108]
  assign _T_3052_data = s2_read ? atomics_data : pstore1_data; // @[DCache.scala 455:108]
  assign _T_3053_opcode = s2_write ? _T_3052_opcode : 3'h4; // @[DCache.scala 455:88]
  assign _T_3053_param = s2_write ? _T_3052_param : 3'h0; // @[DCache.scala 455:88]
  assign _T_3053_size = s2_write ? _T_3052_size : _T_2874_size; // @[DCache.scala 455:88]
  assign _T_3053_source = s2_write ? _T_3052_source : a_source; // @[DCache.scala 455:88]
  assign _T_3053_address = s2_write ? _T_3052_address : s2_req_addr[31:0]; // @[DCache.scala 455:88]
  assign _T_3053_mask = s2_write ? _T_3052_mask : get_mask; // @[DCache.scala 455:88]
  assign _T_3053_data = s2_write ? _T_3052_data : 64'h0; // @[DCache.scala 455:88]
  assign _T_2985_param = {{1'd0}, s2_grow_param}; // @[Edges.scala 323:17 Edges.scala 325:15]
  assign _T_3056 = 2'h1 << a_source; // @[OneHot.scala 52:12]
  assign a_sel = _T_3056[1]; // @[DCache.scala 458:66]
  assign _T_3058 = auto_out_a_ready & tl_out_a_valid; // @[Decoupled.scala 37:37]
  assign _GEN_99 = a_sel | uncachedInFlight_0; // @[DCache.scala 462:18]
  assign _T_3072 = _T_3069 - 9'h1; // @[Edges.scala 230:28]
  assign d_done = d_last & _T_3094; // @[Edges.scala 233:22]
  assign _T_3076 = _T_3067 & ~_T_3072; // @[Edges.scala 234:25]
  assign d_address_inc = {_T_3076, 3'h0}; // @[Edges.scala 269:29]
  assign grantIsVoluntary = auto_out_d_bits_opcode == 3'h6; // @[DCache.scala 490:32]
  assign _T_3089 = blockProbeAfterGrantCount - 3'h1; // @[DCache.scala 494:97]
  assign _T_3096 = cached_grant_wait | reset; // @[DCache.scala 500:13]
  assign _T_3099 = 2'h1 << auto_out_d_bits_source; // @[OneHot.scala 52:12]
  assign d_sel = _T_3099[1]; // @[DCache.scala 508:82]
  assign _T_3103 = d_sel & d_last; // @[DCache.scala 511:17]
  assign _T_3105 = uncachedInFlight_0 | reset; // @[DCache.scala 512:17]
  assign dontCareBits = {tlb_io_resp_paddr[31:3], 3'h0}; // @[DCache.scala 524:53]
  assign _GEN_299 = {{29'd0}, uncachedReqs_0_addr[2:0]}; // @[DCache.scala 525:24]
  assign _T_3110 = dontCareBits | _GEN_299; // @[DCache.scala 525:24]
  assign _T_3112 = release_ack_wait | reset; // @[DCache.scala 530:13]
  assign _GEN_135 = grantIsVoluntary ? 1'h0 : release_ack_wait; // @[DCache.scala 529:36]
  assign _GEN_143 = grantIsUncached ? release_ack_wait : _GEN_135; // @[DCache.scala 507:35]
  assign _GEN_155 = grantIsCached ? release_ack_wait : _GEN_143; // @[DCache.scala 498:26]
  assign _GEN_167 = _T_3094 ? _GEN_155 : release_ack_wait; // @[DCache.scala 497:26]
  assign _T_3114 = auto_out_d_valid & d_first; // @[DCache.scala 536:36]
  assign _T_3115 = _T_3114 & grantIsCached; // @[DCache.scala 536:47]
  assign tl_out__e_valid = _T_3130 ? 1'h0 : _T_3115; // @[DCache.scala 544:51]
  assign _T_3119 = auto_out_e_ready & tl_out__e_valid; // @[Decoupled.scala 37:37]
  assign _T_3121 = _T_3094 & d_first; // @[DCache.scala 538:47]
  assign _T_3122 = _T_3121 & grantIsCached; // @[DCache.scala 538:58]
  assign _T_3123 = _T_3119 == _T_3122; // @[DCache.scala 538:26]
  assign _T_3125 = _T_3123 | reset; // @[DCache.scala 538:9]
  assign _T_3127 = auto_out_d_valid & grantIsRefill; // @[DCache.scala 543:44]
  assign _T_3132 = {s2_vaddr[39:6], 6'h0}; // @[DCache.scala 550:57]
  assign _GEN_300 = {{28'd0}, d_address_inc}; // @[DCache.scala 550:67]
  assign _T_3133 = _T_3132 | _GEN_300; // @[DCache.scala 550:67]
  assign _T_3136 = grantIsCached & d_done; // @[DCache.scala 564:43]
  assign _T_3195 = {s2_write,_T_929,auto_out_d_bits_param}; // @[Cat.scala 30:58]
  assign _T_3204 = 4'hc == _T_3195; // @[Mux.scala 46:19]
  assign _T_3205 = _T_3204 ? 2'h3 : 2'h0; // @[Mux.scala 46:16]
  assign _T_3206 = 4'h4 == _T_3195; // @[Mux.scala 46:19]
  assign _T_3207 = _T_3206 ? 2'h2 : _T_3205; // @[Mux.scala 46:16]
  assign _T_3208 = 4'h0 == _T_3195; // @[Mux.scala 46:19]
  assign _T_3209 = _T_3208 ? 2'h2 : _T_3207; // @[Mux.scala 46:16]
  assign _T_3210 = 4'h1 == _T_3195; // @[Mux.scala 46:19]
  assign _T_3211 = _T_3210 ? 2'h1 : _T_3209; // @[Mux.scala 46:16]
  assign _GEN_170 = auto_out_d_valid ? 1'h0 : _GEN_19; // @[DCache.scala 577:27]
  assign _GEN_171 = auto_out_d_valid | _T_3127; // @[DCache.scala 577:27]
  assign _GEN_172 = auto_out_d_valid ? 1'h0 : 1'h1; // @[DCache.scala 577:27]
  assign _T_3227 = ~block_probe | lrscBackingOff; // @[DCache.scala 588:61]
  assign _T_3228 = auto_out_b_valid & _T_3227; // @[DCache.scala 588:44]
  assign _T_3237 = {io_cpu_req_bits_addr[39:32],auto_out_b_bits_address}; // @[Cat.scala 30:58]
  assign _T_3250 = _T_3247 - 9'h1; // @[Edges.scala 230:28]
  assign c_first = _T_3247 == 9'h0; // @[Edges.scala 231:25]
  assign c_count = _T_3245 & ~_T_3250; // @[Edges.scala 234:25]
  assign releaseRejected = tl_out__c_valid & ~auto_out_c_ready; // @[DCache.scala 598:40]
  assign _T_3261 = {1'h0,c_count}; // @[Cat.scala 30:58]
  assign _T_3262 = {1'h0,s2_release_data_valid}; // @[Cat.scala 30:58]
  assign _GEN_301 = {{1'd0}, s1_release_data_valid}; // @[DCache.scala 601:101]
  assign _T_3264 = _GEN_301 + _T_3262; // @[DCache.scala 601:101]
  assign _T_3265 = releaseRejected ? 2'h0 : _T_3264; // @[DCache.scala 601:52]
  assign _GEN_302 = {{8'd0}, _T_3265}; // @[DCache.scala 601:47]
  assign releaseDataBeat = _T_3261 + _GEN_302; // @[DCache.scala 601:47]
  assign _T_3291 = s2_want_victimize & s2_victim_dirty; // @[DCache.scala 615:24]
  assign _T_3292 = s2_valid & s2_hit_valid; // @[DCache.scala 616:25]
  assign _T_3297 = ~_T_3292 | reset; // @[DCache.scala 616:13]
  assign _T_3300 = {s2_victim_tag,s2_req_addr[11:6]}; // @[Cat.scala 30:58]
  assign res_2_address = {_T_3300, 6'h0}; // @[DCache.scala 618:96]
  assign _GEN_180 = _T_3291 ? 3'h1 : release_state; // @[DCache.scala 615:44]
  assign _T_3305 = releaseDone ? 3'h7 : 3'h3; // @[DCache.scala 629:29]
  assign _T_3307 = releaseDone ? 3'h0 : 3'h5; // @[DCache.scala 633:29]
  assign _GEN_191 = _T_3304 ? s2_report_param : 3'h5; // @[DCache.scala 626:45]
  assign _GEN_197 = _T_3304 ? _T_3305 : _T_3307; // @[DCache.scala 626:45]
  assign _GEN_199 = s2_prb_ack_data ? 3'h2 : _GEN_197; // @[DCache.scala 624:36]
  assign _GEN_202 = s2_prb_ack_data ? 3'h5 : _GEN_191; // @[DCache.scala 624:36]
  assign _GEN_220 = s2_probe ? _GEN_199 : _GEN_180; // @[DCache.scala 620:21]
  assign _GEN_223 = s2_probe ? _GEN_202 : 3'h5; // @[DCache.scala 620:21]
  assign _T_3308 = release_state == 3'h4; // @[DCache.scala 637:25]
  assign _T_3311 = {io_cpu_req_bits_addr[39:32],probe_bits_address}; // @[Cat.scala 30:58]
  assign _GEN_230 = metaArb_io_in_6_ready ? 3'h0 : _GEN_220; // @[DCache.scala 641:37]
  assign _GEN_231 = metaArb_io_in_6_ready | _T_290; // @[DCache.scala 641:37]
  assign _GEN_235 = _T_3308 ? _GEN_230 : _GEN_220; // @[DCache.scala 637:44]
  assign _GEN_237 = releaseDone ? 3'h0 : _GEN_235; // @[DCache.scala 648:26]
  assign _GEN_239 = _T_3312 ? _GEN_237 : _GEN_235; // @[DCache.scala 646:47]
  assign _GEN_243 = _T_3313 ? s2_report_param : _GEN_223; // @[DCache.scala 650:48]
  assign _GEN_252 = _T_3314 ? s2_report_param : _GEN_243; // @[DCache.scala 655:48]
  assign _T_3340 = _T_3238 & c_first; // @[DCache.scala 668:29]
  assign _GEN_260 = _T_3340 | _GEN_167; // @[DCache.scala 668:41]
  assign newCoh_state = _T_3317 ? voluntaryNewCoh_state : probeNewCoh_state; // @[DCache.scala 659:81]
  assign _T_3342 = releaseDataBeat < 10'h8; // @[DCache.scala 676:60]
  assign _T_3345 = {probe_bits_address[11:6], 6'h0}; // @[DCache.scala 679:55]
  assign _T_3347 = {releaseDataBeat[2:0], 3'h0}; // @[DCache.scala 679:117]
  assign _GEN_304 = {{6'd0}, _T_3347}; // @[DCache.scala 679:72]
  assign _T_3352 = release_state == 3'h7; // @[package.scala 14:47]
  assign _T_3362 = metaArb_io_in_4_ready & metaArb_io_in_4_valid; // @[Decoupled.scala 37:37]
  assign _T_3367 = s1_valid | s2_valid; // @[DCache.scala 701:57]
  assign _T_3368 = _T_3367 | cached_grant_wait; // @[DCache.scala 701:94]
  assign _T_3370 = _T_3368 | uncachedInFlight_0; // @[DCache.scala 701:115]
  assign _T_3403 = ~s2_valid_hit_pre_data_ecc | reset; // @[DCache.scala 723:11]
  assign _T_3412 = s2_req_addr[2] ? s2_data_corrected[63:32] : s2_data_corrected[31:0]; // @[AMOALU.scala 39:24]
  assign _T_3415 = a_size == 2'h2; // @[AMOALU.scala 42:26]
  assign _T_3418 = ~s2_req_typ[2] & _T_3412[31]; // @[AMOALU.scala 42:76]
  assign _T_3420 = _T_3418 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  assign _T_3422 = _T_3415 ? _T_3420 : s2_data_corrected[63:32]; // @[AMOALU.scala 42:20]
  assign _T_3423 = {_T_3422,_T_3412}; // @[Cat.scala 30:58]
  assign _T_3427 = s2_req_addr[1] ? _T_3423[31:16] : _T_3423[15:0]; // @[AMOALU.scala 39:24]
  assign _T_3430 = a_size == 2'h1; // @[AMOALU.scala 42:26]
  assign _T_3433 = ~s2_req_typ[2] & _T_3427[15]; // @[AMOALU.scala 42:76]
  assign _T_3435 = _T_3433 ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  assign _T_3437 = _T_3430 ? _T_3435 : _T_3423[63:16]; // @[AMOALU.scala 42:20]
  assign _T_3438 = {_T_3437,_T_3427}; // @[Cat.scala 30:58]
  assign _T_3442 = s2_req_addr[0] ? _T_3438[15:8] : _T_3438[7:0]; // @[AMOALU.scala 39:24]
  assign _T_3444 = _T_752 ? 8'h0 : _T_3442; // @[AMOALU.scala 41:23]
  assign _T_3445 = a_size == 2'h0; // @[AMOALU.scala 42:26]
  assign _T_3446 = _T_3445 | _T_752; // @[AMOALU.scala 42:38]
  assign _T_3448 = ~s2_req_typ[2] & _T_3444[7]; // @[AMOALU.scala 42:76]
  assign _T_3450 = _T_3448 ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  assign _T_3452 = _T_3446 ? _T_3450 : _T_3438[63:8]; // @[AMOALU.scala 42:20]
  assign _T_3453 = {_T_3452,_T_3444}; // @[Cat.scala 30:58]
  assign _GEN_305 = {{63'd0}, s2_sc_fail}; // @[DCache.scala 735:41]
  assign _GEN_290 = _T_3473 | resetting; // @[DCache.scala 759:27]
  assign flushCounterNext = flushCounter + 8'h1; // @[DCache.scala 763:39]
  assign flushDone = flushCounterNext[8:6] == 3'h4; // @[DCache.scala 764:57]
  assign _T_3478 = s2_req_cmd == 5'h5; // @[DCache.scala 766:39]
  assign _T_3479 = s2_valid_masked & _T_3478; // @[DCache.scala 766:25]
  assign _T_3487 = can_acquire_before_release & ~uncachedInFlight_0; // @[DCache.scala 769:56]
  assign _T_3494 = metaArb_io_in_5_ready & metaArb_io_in_5_valid; // @[Decoupled.scala 37:37]
  assign _T_3496 = _T_3494 & ~s1_flush_valid; // @[DCache.scala 774:45]
  assign _T_3498 = _T_3496 & ~s2_flush_valid_pre_tag_ecc; // @[DCache.scala 774:64]
  assign _T_3500 = _T_3498 & _T_357; // @[DCache.scala 774:95]
  assign _T_3505 = {metaArb_io_in_5_bits_idx, 6'h0}; // @[DCache.scala 778:98]
  assign _GEN_295 = resetting ? flushCounterNext : {{1'd0}, flushCounter}; // @[DCache.scala 805:20]
  assign _T_3516 = io_cpu_keep_clock_enabled | metaArb_io_out_valid; // @[DCache.scala 815:31]
  assign _T_3517 = _T_3516 | s1_probe; // @[DCache.scala 816:26]
  assign _T_3518 = _T_3517 | s2_probe; // @[DCache.scala 817:14]
  assign _T_3519 = _T_3518 | s1_valid; // @[DCache.scala 817:26]
  assign _T_3520 = _T_3519 | s2_valid_pre_xcpt; // @[DCache.scala 818:14]
  assign _T_3521 = _T_3520 | pstore1_held; // @[DCache.scala 818:35]
  assign _T_3522 = _T_3521 | pstore2_valid; // @[DCache.scala 819:18]
  assign _T_3524 = _T_3522 | _T_735; // @[DCache.scala 819:35]
  assign _T_3525 = _T_3524 | release_ack_wait; // @[DCache.scala 820:31]
  assign _T_3529 = _T_3525 | ~tlb_io_req_ready; // @[DCache.scala 821:46]
  assign _T_3530 = _T_3529 | cached_grant_wait; // @[DCache.scala 822:23]
  assign _T_3532 = _T_3530 | uncachedInFlight_0; // @[DCache.scala 823:23]
  assign _T_3534 = _T_3532 | _T_1251; // @[DCache.scala 823:54]
  assign auto_out_a_valid = _T_2959 | s2_valid_uncached_pending; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_opcode = s2_uncached ? _T_3053_opcode : 3'h6; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_param = s2_uncached ? _T_3053_param : _T_2985_param; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_size = s2_uncached ? _T_3053_size : 4'h6; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_source = s2_uncached ? _T_3053_source : 1'h0; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_address = s2_uncached ? _T_3053_address : acquire_address[31:0]; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_mask = s2_uncached ? _T_3053_mask : 8'hff; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_data = s2_uncached ? _T_3053_data : 64'h0; // @[LazyModule.scala 173:49]
  assign auto_out_b_ready = _T_3232 & ~s2_valid; // @[LazyModule.scala 173:49]
  assign auto_out_c_valid = _T_3313 | _GEN_238; // @[LazyModule.scala 173:49]
  assign auto_out_c_bits_opcode = _T_3317 ? 3'h7 : _GEN_251; // @[LazyModule.scala 173:49]
  assign auto_out_c_bits_param = _T_3317 ? s2_shrink_param : _GEN_252; // @[LazyModule.scala 173:49]
  assign auto_out_c_bits_size = _T_3317 ? 4'h6 : probe_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_c_bits_source = probe_bits_source; // @[LazyModule.scala 173:49]
  assign auto_out_c_bits_address = probe_bits_address; // @[LazyModule.scala 173:49]
  assign auto_out_c_bits_data = {_T_1026,_T_1023}; // @[LazyModule.scala 173:49]
  assign auto_out_d_ready = _T_3219 ? 1'h0 : _GEN_169; // @[LazyModule.scala 173:49]
  assign auto_out_e_valid = _T_3130 ? 1'h0 : _T_3115; // @[LazyModule.scala 173:49]
  assign auto_out_e_bits_sink = auto_out_d_bits_sink; // @[LazyModule.scala 173:49]
  assign io_cpu_req_ready = _T_3219 ? _GEN_170 : _GEN_19; // @[DCache.scala 159:20 DCache.scala 173:64 DCache.scala 181:53 DCache.scala 192:98 DCache.scala 578:24]
  assign io_cpu_s2_nack = _T_3479 ? ~flushed : _T_1200; // @[DCache.scala 300:18 DCache.scala 767:20]
  assign io_cpu_resp_valid = doUncachedResp | s2_valid_hit_pre_data_ecc; // @[DCache.scala 692:21 DCache.scala 724:23]
  assign io_cpu_resp_bits_tag = s2_req_tag; // @[DCache.scala 693:20]
  assign io_cpu_resp_bits_typ = s2_req_typ; // @[DCache.scala 693:20]
  assign io_cpu_resp_bits_data = _T_3453 | _GEN_305; // @[DCache.scala 693:20 DCache.scala 735:25]
  assign io_cpu_resp_bits_replay = doUncachedResp; // @[DCache.scala 695:27 DCache.scala 725:29]
  assign io_cpu_resp_bits_has_data = _T_753 | _T_770; // @[DCache.scala 694:29]
  assign io_cpu_resp_bits_data_word_bypass = {_T_3422,_T_3412}; // @[DCache.scala 736:37]
  assign io_cpu_replay_next = _T_3094 & grantIsUncachedData; // @[DCache.scala 719:22]
  assign io_cpu_s2_xcpt_ma_ld = _T_3374 & _T_3376_ma_ld; // @[DCache.scala 705:18]
  assign io_cpu_s2_xcpt_ma_st = _T_3374 & _T_3376_ma_st; // @[DCache.scala 705:18]
  assign io_cpu_s2_xcpt_pf_ld = _T_3374 & _T_3376_pf_ld; // @[DCache.scala 705:18]
  assign io_cpu_s2_xcpt_pf_st = _T_3374 & _T_3376_pf_st; // @[DCache.scala 705:18]
  assign io_cpu_s2_xcpt_ae_ld = _T_3374 & _T_3376_ae_ld; // @[DCache.scala 705:18]
  assign io_cpu_s2_xcpt_ae_st = _T_3374 & _T_3376_ae_st; // @[DCache.scala 705:18]
  assign io_cpu_ordered = ~_T_3370; // @[DCache.scala 701:18]
  assign io_cpu_perf_grant = d_last & _T_3094; // @[DCache.scala 829:21]
  assign io_cpu_clock_enabled = clock_en_reg; // @[DCache.scala 89:24]
  assign io_ptw_req_valid = tlb_io_ptw_req_valid; // @[DCache.scala 185:10]
  assign io_ptw_req_bits_bits_addr = tlb_io_ptw_req_bits_bits_addr; // @[DCache.scala 185:10]
  assign metaArb_io_in_0_valid = resetting; // @[DCache.scala 800:26]
  assign metaArb_io_in_0_bits_addr = metaArb_io_in_5_bits_addr; // @[DCache.scala 801:25]
  assign metaArb_io_in_0_bits_idx = metaArb_io_in_5_bits_idx; // @[DCache.scala 801:25]
  assign metaArb_io_in_0_bits_data = {2'h0,s2_req_addr[31:12]}; // @[DCache.scala 801:25 DCache.scala 804:30]
  assign metaArb_io_in_2_valid = _T_1201 | _T_1234; // @[DCache.scala 317:26]
  assign metaArb_io_in_2_bits_addr = {io_cpu_req_bits_addr[39:12],s2_vaddr[11:0]}; // @[DCache.scala 321:30]
  assign metaArb_io_in_2_bits_idx = s2_vaddr[11:6]; // @[DCache.scala 320:29]
  assign metaArb_io_in_2_bits_way_en = s2_hit_valid ? s2_hit_way : _T_1061; // @[DCache.scala 319:32]
  assign metaArb_io_in_2_bits_data = {_T_1244_state,s2_req_addr[31:12]}; // @[DCache.scala 322:30]
  assign metaArb_io_in_3_valid = _T_3136 & ~auto_out_d_bits_denied; // @[DCache.scala 564:26]
  assign metaArb_io_in_3_bits_addr = {io_cpu_req_bits_addr[39:12],s2_vaddr[11:0]}; // @[DCache.scala 568:30]
  assign metaArb_io_in_3_bits_idx = s2_vaddr[11:6]; // @[DCache.scala 567:29]
  assign metaArb_io_in_3_bits_way_en = s2_hit_valid ? s2_hit_way : _T_1061; // @[DCache.scala 566:32]
  assign metaArb_io_in_3_bits_data = {_T_3211,s2_req_addr[31:12]}; // @[DCache.scala 569:30]
  assign metaArb_io_in_4_valid = _T_3316 | _T_3352; // @[DCache.scala 683:26]
  assign metaArb_io_in_4_bits_addr = {io_cpu_req_bits_addr[39:12],probe_bits_address[11:0]}; // @[DCache.scala 687:30]
  assign metaArb_io_in_4_bits_idx = probe_bits_address[11:6]; // @[DCache.scala 686:29]
  assign metaArb_io_in_4_bits_way_en = _T_3317 ? s2_victim_way : s2_probe_way; // @[DCache.scala 685:32]
  assign metaArb_io_in_4_bits_data = {newCoh_state,probe_bits_address[31:12]}; // @[DCache.scala 688:30]
  assign metaArb_io_in_5_valid = flushing; // @[DCache.scala 775:26]
  assign metaArb_io_in_5_bits_addr = {io_cpu_req_bits_addr[39:12],_T_3505}; // @[DCache.scala 778:30]
  assign metaArb_io_in_5_bits_idx = flushCounter[5:0]; // @[DCache.scala 777:29]
  assign metaArb_io_in_5_bits_way_en = metaArb_io_in_4_bits_way_en; // @[DCache.scala 779:32]
  assign metaArb_io_in_5_bits_data = metaArb_io_in_4_bits_data; // @[DCache.scala 780:30]
  assign metaArb_io_in_6_valid = _T_3308 | _T_3228; // @[DCache.scala 588:26 DCache.scala 638:30]
  assign metaArb_io_in_6_bits_addr = _T_3308 ? _T_3311 : _T_3237; // @[DCache.scala 592:30 DCache.scala 640:34]
  assign metaArb_io_in_6_bits_idx = _T_3308 ? probe_bits_address[11:6] : auto_out_b_bits_address[11:6]; // @[DCache.scala 591:29 DCache.scala 639:33]
  assign metaArb_io_in_6_bits_way_en = metaArb_io_in_4_bits_way_en; // @[DCache.scala 593:32]
  assign metaArb_io_in_6_bits_data = metaArb_io_in_4_bits_data; // @[DCache.scala 594:30]
  assign metaArb_io_in_7_valid = io_cpu_req_valid; // @[DCache.scala 175:26]
  assign metaArb_io_in_7_bits_addr = io_cpu_req_bits_addr; // @[DCache.scala 178:30]
  assign metaArb_io_in_7_bits_idx = io_cpu_req_bits_addr[11:6]; // @[DCache.scala 177:29]
  assign metaArb_io_in_7_bits_way_en = metaArb_io_in_4_bits_way_en; // @[DCache.scala 179:32]
  assign metaArb_io_in_7_bits_data = metaArb_io_in_4_bits_data; // @[DCache.scala 180:30]
  assign metaArb_io_out_ready = clock_en_reg; // @[DCache.scala 114:24]
  assign data_clock = gated_clock;
  assign data_io_req_valid = dataArb_io_out_valid; // @[DCache.scala 111:15]
  assign data_io_req_bits_addr = dataArb_io_out_bits_addr; // @[DCache.scala 111:15]
  assign data_io_req_bits_write = dataArb_io_out_bits_write; // @[DCache.scala 111:15]
  assign data_io_req_bits_wdata = {_T_284,_T_281}; // @[DCache.scala 111:15 DCache.scala 112:26]
  assign data_io_req_bits_eccMask = dataArb_io_out_bits_eccMask; // @[DCache.scala 111:15]
  assign data_io_req_bits_way_en = dataArb_io_out_bits_way_en; // @[DCache.scala 111:15]
  assign dataArb_io_in_0_valid = pstore_drain_structural | _T_1460; // @[DCache.scala 403:26]
  assign dataArb_io_in_0_bits_addr = _T_1560[11:0]; // @[DCache.scala 405:30]
  assign dataArb_io_in_0_bits_write = pstore_drain_structural | _T_1460; // @[DCache.scala 404:31]
  assign dataArb_io_in_0_bits_wdata = pstore2_valid ? pstore2_storegen_data : pstore1_data; // @[DCache.scala 407:31]
  assign dataArb_io_in_0_bits_eccMask = {_T_1587,_T_1584}; // @[DCache.scala 410:33]
  assign dataArb_io_in_0_bits_way_en = pstore2_valid ? pstore2_way : pstore1_way; // @[DCache.scala 406:32]
  assign dataArb_io_in_1_valid = _T_3219 ? _GEN_171 : _T_3127; // @[DCache.scala 543:26 DCache.scala 579:30]
  assign dataArb_io_in_1_bits_addr = _T_3133[11:0]; // @[DCache.scala 550:32]
  assign dataArb_io_in_1_bits_write = _T_3219 ? _GEN_172 : 1'h1; // @[DCache.scala 549:33 DCache.scala 580:35]
  assign dataArb_io_in_1_bits_wdata = auto_out_d_bits_data; // @[DCache.scala 110:43 DCache.scala 552:33]
  assign dataArb_io_in_1_bits_eccMask = 8'hff; // @[DCache.scala 555:35]
  assign dataArb_io_in_1_bits_way_en = s2_hit_valid ? s2_hit_way : _T_1061; // @[DCache.scala 551:34]
  assign dataArb_io_in_2_valid = inWriteback & _T_3342; // @[DCache.scala 676:26]
  assign dataArb_io_in_2_bits_addr = _T_3345 | _GEN_304; // @[DCache.scala 677:25 DCache.scala 679:30]
  assign dataArb_io_in_2_bits_wdata = dataArb_io_in_1_bits_wdata; // @[DCache.scala 110:43 DCache.scala 677:25]
  assign dataArb_io_in_2_bits_eccMask = dataArb_io_in_1_bits_eccMask; // @[DCache.scala 677:25]
  assign dataArb_io_in_3_valid = io_cpu_req_valid & res; // @[DCache.scala 167:26]
  assign dataArb_io_in_3_bits_addr = io_cpu_req_bits_addr[11:0]; // @[DCache.scala 168:25 DCache.scala 170:30]
  assign dataArb_io_in_3_bits_wdata = dataArb_io_in_1_bits_wdata; // @[DCache.scala 110:43 DCache.scala 168:25]
  assign dataArb_io_in_3_bits_eccMask = dataArb_io_in_1_bits_eccMask; // @[DCache.scala 168:25]
  assign tlb_clock = gated_clock;
  assign tlb_reset = reset;
  assign tlb_io_req_valid = s1_valid_masked & s1_readwrite; // @[DCache.scala 187:20]
  assign tlb_io_req_bits_vaddr = s1_req_addr; // @[DCache.scala 189:25]
  assign tlb_io_req_bits_passthrough = s1_req_phys; // @[DCache.scala 188:31]
  assign tlb_io_req_bits_size = s1_req_typ[1:0]; // @[DCache.scala 190:24]
  assign tlb_io_req_bits_cmd = s1_req_cmd; // @[DCache.scala 191:23]
  assign tlb_io_sfence_valid = s1_valid_masked & s1_sfence; // @[DCache.scala 195:23]
  assign tlb_io_sfence_bits_rs1 = s1_req_typ[0]; // @[DCache.scala 196:26]
  assign tlb_io_sfence_bits_rs2 = s1_req_typ[1]; // @[DCache.scala 197:26]
  assign tlb_io_sfence_bits_addr = s1_req_addr[38:0]; // @[DCache.scala 199:27]
  assign tlb_io_ptw_req_ready = io_ptw_req_ready; // @[DCache.scala 185:10]
  assign tlb_io_ptw_resp_valid = io_ptw_resp_valid; // @[DCache.scala 185:10]
  assign tlb_io_ptw_resp_bits_ae = io_ptw_resp_bits_ae; // @[DCache.scala 185:10]
  assign tlb_io_ptw_resp_bits_pte_ppn = io_ptw_resp_bits_pte_ppn; // @[DCache.scala 185:10]
  assign tlb_io_ptw_resp_bits_pte_d = io_ptw_resp_bits_pte_d; // @[DCache.scala 185:10]
  assign tlb_io_ptw_resp_bits_pte_a = io_ptw_resp_bits_pte_a; // @[DCache.scala 185:10]
  assign tlb_io_ptw_resp_bits_pte_g = io_ptw_resp_bits_pte_g; // @[DCache.scala 185:10]
  assign tlb_io_ptw_resp_bits_pte_u = io_ptw_resp_bits_pte_u; // @[DCache.scala 185:10]
  assign tlb_io_ptw_resp_bits_pte_x = io_ptw_resp_bits_pte_x; // @[DCache.scala 185:10]
  assign tlb_io_ptw_resp_bits_pte_w = io_ptw_resp_bits_pte_w; // @[DCache.scala 185:10]
  assign tlb_io_ptw_resp_bits_pte_r = io_ptw_resp_bits_pte_r; // @[DCache.scala 185:10]
  assign tlb_io_ptw_resp_bits_pte_v = io_ptw_resp_bits_pte_v; // @[DCache.scala 185:10]
  assign tlb_io_ptw_resp_bits_level = io_ptw_resp_bits_level; // @[DCache.scala 185:10]
  assign tlb_io_ptw_resp_bits_homogeneous = io_ptw_resp_bits_homogeneous; // @[DCache.scala 185:10]
  assign tlb_io_ptw_ptbr_mode = io_ptw_ptbr_mode; // @[DCache.scala 185:10]
  assign tlb_io_ptw_status_dprv = io_ptw_status_dprv; // @[DCache.scala 185:10]
  assign tlb_io_ptw_status_mxr = io_ptw_status_mxr; // @[DCache.scala 185:10]
  assign tlb_io_ptw_status_sum = io_ptw_status_sum; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_0_addr = io_ptw_pmp_0_addr; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_0_mask = io_ptw_pmp_0_mask; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_1_addr = io_ptw_pmp_1_addr; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_1_mask = io_ptw_pmp_1_mask; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_2_addr = io_ptw_pmp_2_addr; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_2_mask = io_ptw_pmp_2_mask; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_3_addr = io_ptw_pmp_3_addr; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_3_mask = io_ptw_pmp_3_mask; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_4_addr = io_ptw_pmp_4_addr; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_4_mask = io_ptw_pmp_4_mask; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_5_addr = io_ptw_pmp_5_addr; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_5_mask = io_ptw_pmp_5_mask; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_6_addr = io_ptw_pmp_6_addr; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_6_mask = io_ptw_pmp_6_mask; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_7_addr = io_ptw_pmp_7_addr; // @[DCache.scala 185:10]
  assign tlb_io_ptw_pmp_7_mask = io_ptw_pmp_7_mask; // @[DCache.scala 185:10]
  assign tlb_io_ptw_vpoffset_bits_value = io_ptw_vpoffset_bits_value; // @[DCache.scala 185:10]
  assign amoalu_io_mask = pstore1_mask; // @[DCache.scala 744:20]
  assign amoalu_io_cmd = pstore1_cmd; // @[DCache.scala 745:19]
  assign amoalu_io_lhs = {_T_1026,_T_1023}; // @[DCache.scala 746:19]
  assign amoalu_io_rhs = pstore1_data; // @[DCache.scala 747:19]
  assign _GEN_308 = _T_3094 & grantIsCached; // @[DCache.scala 500:13]
  assign _GEN_311 = _T_3094 & ~grantIsCached; // @[DCache.scala 512:17]
  assign _GEN_312 = _GEN_311 & grantIsUncached; // @[DCache.scala 512:17]
  assign _GEN_313 = _GEN_312 & _T_3103; // @[DCache.scala 512:17]
  assign _GEN_321 = _GEN_311 & ~grantIsUncached; // @[DCache.scala 530:13]
  assign _GEN_322 = _GEN_321 & grantIsVoluntary; // @[DCache.scala 530:13]
  assign DCache_cov_read_addr = DCache_state;
  assign DCache_cov_read_data = DCache_cov[DCache_cov_read_addr]; // @[Coverage map for DCache]
  assign DCache_cov_write_data = 1'h1;
  assign DCache_cov_write_addr = DCache_state;
  assign DCache_cov_write_mask = 1'h1;
  assign DCache_cov_write_en = 1'h1;
  assign mux_cond_0 = s1_req_addr[1];
  assign mux_cond_1 = s2_req_addr[0];
  assign mux_cond_2 = s2_req_addr[2];
  assign mux_cond_3 = s1_req_addr[2];
  assign mux_cond_4 = s2_req_addr[1];
  assign mux_cond_5 = s1_req_addr[0];
  assign pstore1_held_shl = {pstore1_held, 18'h0};
  assign pstore1_held_pad = {1'h0,pstore1_held_shl};
  assign s2_valid_pre_xcpt_shl = {s2_valid_pre_xcpt, 15'h0};
  assign s2_valid_pre_xcpt_pad = {4'h0,s2_valid_pre_xcpt_shl};
  assign s2_release_data_valid_shl = {s2_release_data_valid, 7'h0};
  assign s2_release_data_valid_pad = {12'h0,s2_release_data_valid_shl};
  assign s2_flush_valid_pre_tag_ecc_shl = {s2_flush_valid_pre_tag_ecc, 15'h0};
  assign s2_flush_valid_pre_tag_ecc_pad = {4'h0,s2_flush_valid_pre_tag_ecc_shl};
  assign s2_hit_way_shl = {s2_hit_way, 11'h0};
  assign s2_hit_way_pad = {5'h0,s2_hit_way_shl};
  assign _T_1060_shl = {_T_1060, 3'h0};
  assign _T_1060_pad = {15'h0,_T_1060_shl};
  assign s2_hit_state_state_shl = {s2_hit_state_state, 11'h0};
  assign s2_hit_state_state_pad = {7'h0,s2_hit_state_state_shl};
  assign pstore2_valid_shl = {pstore2_valid, 18'h0};
  assign pstore2_valid_pad = {1'h0,pstore2_valid_shl};
  assign uncachedInFlight_0_shl = {uncachedInFlight_0, 15'h0};
  assign uncachedInFlight_0_pad = {4'h0,uncachedInFlight_0_shl};
  assign s2_probe_shl = {s2_probe, 6'h0};
  assign s2_probe_pad = {13'h0,s2_probe_shl};
  assign resetting_shl = {resetting, 12'h0};
  assign resetting_pad = {7'h0,resetting_shl};
  assign s2_probe_way_shl = {s2_probe_way, 1'h0};
  assign s2_probe_way_pad = {15'h0,s2_probe_way_shl};
  assign s1_valid_shl = {s1_valid, 12'h0};
  assign s1_valid_pad = {7'h0,s1_valid_shl};
  assign grantInProgress_shl = {grantInProgress, 18'h0};
  assign grantInProgress_pad = {1'h0,grantInProgress_shl};
  assign s2_req_typ_shl = {s2_req_typ, 8'h0};
  assign s2_req_typ_pad = {9'h0,s2_req_typ_shl};
  assign s2_probe_state_state_shl = s2_probe_state_state;
  assign s2_probe_state_state_pad = {18'h0,s2_probe_state_state_shl};
  assign cached_grant_wait_shl = {cached_grant_wait, 3'h0};
  assign cached_grant_wait_pad = {16'h0,cached_grant_wait_shl};
  assign flushed_shl = {flushed, 12'h0};
  assign flushed_pad = {7'h0,flushed_shl};
  assign release_ack_wait_shl = {release_ack_wait, 5'h0};
  assign release_ack_wait_pad = {14'h0,release_ack_wait_shl};
  assign s2_uncached_shl = {s2_uncached, 15'h0};
  assign s2_uncached_pad = {4'h0,s2_uncached_shl};
  assign release_state_shl = {release_state, 17'h0};
  assign release_state_pad = release_state_shl;
  assign s1_flush_valid_shl = {s1_flush_valid, 16'h0};
  assign s1_flush_valid_pad = {3'h0,s1_flush_valid_shl};
  assign blockUncachedGrant_shl = {blockUncachedGrant, 4'h0};
  assign blockUncachedGrant_pad = {15'h0,blockUncachedGrant_shl};
  assign _T_1068_state_shl = _T_1068_state;
  assign _T_1068_state_pad = {18'h0,_T_1068_state_shl};
  assign _T_738_shl = {_T_738, 1'h0};
  assign _T_738_pad = {18'h0,_T_738_shl};
  assign probe_bits_param_shl = {probe_bits_param, 14'h0};
  assign probe_bits_param_pad = {4'h0,probe_bits_param_shl};
  assign s1_probe_shl = {s1_probe, 4'h0};
  assign s1_probe_pad = {15'h0,s1_probe_shl};
  assign pstore1_rmw_shl = {pstore1_rmw, 6'h0};
  assign pstore1_rmw_pad = {13'h0,pstore1_rmw_shl};
  assign s1_req_typ_shl = {s1_req_typ, 14'h0};
  assign s1_req_typ_pad = {3'h0,s1_req_typ_shl};
  assign mux_cond_0_shl = {mux_cond_0, 11'h0};
  assign mux_cond_0_pad = {8'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 10'h0};
  assign mux_cond_1_pad = {9'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 1'h0};
  assign mux_cond_2_pad = {18'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 12'h0};
  assign mux_cond_3_pad = {7'h0,mux_cond_3_shl};
  assign mux_cond_4_shl = {mux_cond_4, 17'h0};
  assign mux_cond_4_pad = {2'h0,mux_cond_4_shl};
  assign mux_cond_5_shl = {mux_cond_5, 2'h0};
  assign mux_cond_5_pad = {17'h0,mux_cond_5_shl};
  assign DCache_xor15 = pstore1_held_pad ^ s2_valid_pre_xcpt_pad;
  assign DCache_xor16 = s2_release_data_valid_pad ^ s2_flush_valid_pre_tag_ecc_pad;
  assign DCache_xor7 = DCache_xor15 ^ DCache_xor16;
  assign DCache_xor17 = s2_hit_way_pad ^ _T_1060_pad;
  assign DCache_xor18 = s2_hit_state_state_pad ^ pstore2_valid_pad;
  assign DCache_xor8 = DCache_xor17 ^ DCache_xor18;
  assign DCache_xor3 = DCache_xor7 ^ DCache_xor8;
  assign DCache_xor19 = uncachedInFlight_0_pad ^ s2_probe_pad;
  assign DCache_xor20 = resetting_pad ^ s2_probe_way_pad;
  assign DCache_xor9 = DCache_xor19 ^ DCache_xor20;
  assign DCache_xor21 = s1_valid_pad ^ grantInProgress_pad;
  assign DCache_xor46 = s2_probe_state_state_pad ^ cached_grant_wait_pad;
  assign DCache_xor22 = s2_req_typ_pad ^ DCache_xor46;
  assign DCache_xor10 = DCache_xor21 ^ DCache_xor22;
  assign DCache_xor4 = DCache_xor9 ^ DCache_xor10;
  assign DCache_xor1 = DCache_xor3 ^ DCache_xor4;
  assign DCache_xor23 = flushed_pad ^ release_ack_wait_pad;
  assign DCache_xor24 = s2_uncached_pad ^ release_state_pad;
  assign DCache_xor11 = DCache_xor23 ^ DCache_xor24;
  assign DCache_xor25 = s1_flush_valid_pad ^ blockUncachedGrant_pad;
  assign DCache_xor54 = _T_738_pad ^ probe_bits_param_pad;
  assign DCache_xor26 = _T_1068_state_pad ^ DCache_xor54;
  assign DCache_xor12 = DCache_xor25 ^ DCache_xor26;
  assign DCache_xor5 = DCache_xor11 ^ DCache_xor12;
  assign DCache_xor27 = s1_probe_pad ^ pstore1_rmw_pad;
  assign DCache_xor28 = s1_req_typ_pad ^ mux_cond_0_pad;
  assign DCache_xor13 = DCache_xor27 ^ DCache_xor28;
  assign DCache_xor29 = mux_cond_1_pad ^ mux_cond_2_pad;
  assign DCache_xor62 = mux_cond_4_pad ^ mux_cond_5_pad;
  assign DCache_xor30 = mux_cond_3_pad ^ DCache_xor62;
  assign DCache_xor14 = DCache_xor29 ^ DCache_xor30;
  assign DCache_xor6 = DCache_xor13 ^ DCache_xor14;
  assign DCache_xor2 = DCache_xor5 ^ DCache_xor6;
  assign DCache_xor0 = DCache_xor1 ^ DCache_xor2;
  assign dataArb_sum = DCache_covSum + dataArb_io_covSum;
  assign amoalu_sum = dataArb_sum + amoalu_io_covSum;
  assign data_sum = amoalu_sum + data_io_covSum;
  assign metaArb_sum = data_sum + metaArb_io_covSum;
  assign tlb_sum = metaArb_sum + tlb_io_covSum;
  assign io_covSum = tlb_sum;
  assign stopEn0 = ~_T_471;
  assign stopEn1 = ~_T_471;
  assign stopEn2 = ~_T_1441;
  assign stopEn3 = _GEN_308 & ~_T_3096;
  assign stopEn4 = _GEN_313 & ~_T_3105;
  assign stopEn5 = _GEN_322 & ~_T_3112;
  assign stopEn6 = ~_T_3125;
  assign stopEn7 = _T_3291 & ~_T_3297;
  assign stopEn8 = doUncachedResp & ~_T_3403;
  assign amoalu_metaAssert_wire = amoalu_metaAssert;
  assign dataArb_metaAssert_wire = dataArb_metaAssert;
  assign data_metaAssert_wire = data_metaAssert;
  assign tlb_metaAssert_wire = tlb_metaAssert;
  assign metaArb_metaAssert_wire = metaArb_metaAssert;
  assign DCache_or8 = stopEn1 | stopEn2;
  assign DCache_or3 = stopEn0 | DCache_or8;
  assign DCache_or9 = stopEn3 | stopEn4;
  assign DCache_or10 = stopEn5 | stopEn6;
  assign DCache_or4 = DCache_or9 | DCache_or10;
  assign DCache_or1 = DCache_or3 | DCache_or4;
  assign DCache_or12 = stopEn8 | dataArb_metaAssert_wire;
  assign DCache_or5 = stopEn7 | DCache_or12;
  assign DCache_or13 = tlb_metaAssert_wire | amoalu_metaAssert_wire;
  assign DCache_or14 = data_metaAssert_wire | metaArb_metaAssert_wire;
  assign DCache_or6 = DCache_or13 | DCache_or14;
  assign DCache_or2 = DCache_or5 | DCache_or6;
  assign DCache_or0 = DCache_or1 | DCache_or2;
  assign metaAssert = DCache_or0;
  assign data_metaReset = metaReset | data_halt;
  assign tlb_metaReset = metaReset | tlb_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_0[initvar] = _RAND_0[21:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tag_array_0_s1_meta_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  tag_array_0_s1_meta_addr_pipe_0 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_1[initvar] = _RAND_3[21:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  tag_array_1_s1_meta_en_pipe_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  tag_array_1_s1_meta_addr_pipe_0 = _RAND_5[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_2[initvar] = _RAND_6[21:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  tag_array_2_s1_meta_en_pipe_0 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  tag_array_2_s1_meta_addr_pipe_0 = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_3[initvar] = _RAND_9[21:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  tag_array_3_s1_meta_en_pipe_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  tag_array_3_s1_meta_addr_pipe_0 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  clock_en_reg = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  lfsr = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  blockUncachedGrant = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  s1_valid = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_3069 = _RAND_16[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  s1_probe = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  s2_probe = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  release_state = _RAND_19[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  grantInProgress = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  blockProbeAfterGrantCount = _RAND_21[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  lrscCount = _RAND_22[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  s2_valid_pre_xcpt = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  probe_bits_param = _RAND_24[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  probe_bits_size = _RAND_25[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  probe_bits_source = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  probe_bits_address = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  s2_probe_state_state = _RAND_28[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_3247 = _RAND_29[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  s2_release_data_valid = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  s1_req_cmd = _RAND_31[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_738 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  s2_req_cmd = _RAND_33[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  s2_hit_state_state = _RAND_34[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {2{`RANDOM}};
  lrscAddr = _RAND_35[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {2{`RANDOM}};
  s2_req_addr = _RAND_36[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  pstore1_held = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {2{`RANDOM}};
  pstore1_addr = _RAND_38[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{`RANDOM}};
  s1_req_addr = _RAND_39[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  pstore1_mask = _RAND_40[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  s1_req_typ = _RAND_41[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  pstore2_valid = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {2{`RANDOM}};
  pstore2_addr = _RAND_43[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  mask = _RAND_44[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  s1_req_tag = _RAND_45[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  s1_req_phys = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  s1_flush_valid = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  cached_grant_wait = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  release_ack_wait = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  uncachedInFlight_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {2{`RANDOM}};
  uncachedReqs_0_addr = _RAND_51[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  uncachedReqs_0_tag = _RAND_52[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  uncachedReqs_0_typ = _RAND_53[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  s2_hit_way = _RAND_54[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_1060 = _RAND_55[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  s2_probe_way = _RAND_56[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  s2_req_tag = _RAND_57[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  s2_req_typ = _RAND_58[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  s2_uncached = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {2{`RANDOM}};
  _T_746 = _RAND_60[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  s2_flush_valid_pre_tag_ecc = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {2{`RANDOM}};
  s2_data = _RAND_62[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  s2_victim_tag = _RAND_63[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_1068_state = _RAND_64[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  pstore1_cmd = _RAND_65[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {2{`RANDOM}};
  pstore1_data = _RAND_66[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  pstore1_way = _RAND_67[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  pstore1_rmw = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  pstore2_way = _RAND_69[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_1487 = _RAND_70[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_1493 = _RAND_71[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_1499 = _RAND_72[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_1505 = _RAND_73[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_1511 = _RAND_74[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_1517 = _RAND_75[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_1523 = _RAND_76[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_1529 = _RAND_77[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  s1_release_data_valid = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_3374 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_3376_pf_ld = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_3376_pf_st = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_3376_ae_ld = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_3376_ae_st = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_3376_ma_ld = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_3376_ma_st = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  doUncachedResp = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  resetting = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_3473 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  flushed = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  flushing = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  flushCounter = _RAND_91[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  DCache_state = _RAND_92[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    DCache_cov[initvar] = _RAND_93[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  DCache_covSum = _RAND_94[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge gated_clock) begin
    if(tag_array_0__T_567_en & tag_array_0__T_567_mask) begin
      tag_array_0[tag_array_0__T_567_addr] <= tag_array_0__T_567_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      tag_array_0_s1_meta_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_0_s1_meta_en_pipe_0 <= metaArb_io_out_valid & ~metaArb_io_out_bits_write;
    end
    if (metaReset) begin
      tag_array_0_s1_meta_addr_pipe_0 <= 6'h0;
    end else if (metaArb_io_out_valid & ~metaArb_io_out_bits_write) begin
      tag_array_0_s1_meta_addr_pipe_0 <= metaArb_io_out_bits_idx;
    end
    if(tag_array_1__T_567_en & tag_array_1__T_567_mask) begin
      tag_array_1[tag_array_1__T_567_addr] <= tag_array_1__T_567_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      tag_array_1_s1_meta_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_1_s1_meta_en_pipe_0 <= metaArb_io_out_valid & ~metaArb_io_out_bits_write;
    end
    if (metaReset) begin
      tag_array_1_s1_meta_addr_pipe_0 <= 6'h0;
    end else if (metaArb_io_out_valid & ~metaArb_io_out_bits_write) begin
      tag_array_1_s1_meta_addr_pipe_0 <= metaArb_io_out_bits_idx;
    end
    if(tag_array_2__T_567_en & tag_array_2__T_567_mask) begin
      tag_array_2[tag_array_2__T_567_addr] <= tag_array_2__T_567_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      tag_array_2_s1_meta_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_2_s1_meta_en_pipe_0 <= metaArb_io_out_valid & ~metaArb_io_out_bits_write;
    end
    if (metaReset) begin
      tag_array_2_s1_meta_addr_pipe_0 <= 6'h0;
    end else if (metaArb_io_out_valid & ~metaArb_io_out_bits_write) begin
      tag_array_2_s1_meta_addr_pipe_0 <= metaArb_io_out_bits_idx;
    end
    if(tag_array_3__T_567_en & tag_array_3__T_567_mask) begin
      tag_array_3[tag_array_3__T_567_addr] <= tag_array_3__T_567_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      tag_array_3_s1_meta_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_3_s1_meta_en_pipe_0 <= metaArb_io_out_valid & ~metaArb_io_out_bits_write;
    end
    if (metaReset) begin
      tag_array_3_s1_meta_addr_pipe_0 <= 6'h0;
    end else if (metaArb_io_out_valid & ~metaArb_io_out_bits_write) begin
      tag_array_3_s1_meta_addr_pipe_0 <= metaArb_io_out_bits_idx;
    end
    if (metaReset) begin
      clock_en_reg <= 1'h0;
    end else begin
      clock_en_reg <= _T_3534 | _T_3224;
    end
    if (metaReset) begin
      lfsr <= 16'h0;
    end else if (reset) begin
      lfsr <= 16'h1;
    end else if (_GEN_159) begin
      lfsr <= _T_257;
    end
    if (metaReset) begin
      blockUncachedGrant <= 1'h0;
    end else if (_T_3219) begin
      if (auto_out_d_valid) begin
        blockUncachedGrant <= ~dataArb_io_in_1_ready;
      end else begin
        blockUncachedGrant <= dataArb_io_out_valid;
      end
    end else begin
      blockUncachedGrant <= dataArb_io_out_valid;
    end
    if (metaReset) begin
      s1_valid <= 1'h0;
    end else if (reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= _T_288;
    end
    if (metaReset) begin
      _T_3069 <= 9'h0;
    end else if (reset) begin
      _T_3069 <= 9'h0;
    end else if (_T_3094) begin
      if (d_first) begin
        if (auto_out_d_bits_opcode[0]) begin
          _T_3069 <= _T_3065;
        end else begin
          _T_3069 <= 9'h0;
        end
      end else begin
        _T_3069 <= _T_3072;
      end
    end
    if (metaReset) begin
      s1_probe <= 1'h0;
    end else if (reset) begin
      s1_probe <= 1'h0;
    end else if (_T_3308) begin
      s1_probe <= _GEN_231;
    end else begin
      s1_probe <= _T_290;
    end
    if (metaReset) begin
      s2_probe <= 1'h0;
    end else if (reset) begin
      s2_probe <= 1'h0;
    end else begin
      s2_probe <= s1_probe;
    end
    if (metaReset) begin
      release_state <= 3'h0;
    end else if (reset) begin
      release_state <= 3'h0;
    end else if (_T_3362) begin
      release_state <= 3'h0;
    end else if (_T_3317) begin
      if (releaseDone) begin
        release_state <= 3'h6;
      end else if (_T_3314) begin
        if (releaseDone) begin
          release_state <= 3'h7;
        end else if (_T_3313) begin
          if (releaseDone) begin
            release_state <= 3'h7;
          end else if (_T_3312) begin
            if (releaseDone) begin
              release_state <= 3'h0;
            end else if (_T_3308) begin
              if (metaArb_io_in_6_ready) begin
                release_state <= 3'h0;
              end else if (s2_probe) begin
                if (s2_prb_ack_data) begin
                  release_state <= 3'h2;
                end else if (_T_3304) begin
                  if (releaseDone) begin
                    release_state <= 3'h7;
                  end else begin
                    release_state <= 3'h3;
                  end
                end else if (releaseDone) begin
                  release_state <= 3'h0;
                end else begin
                  release_state <= 3'h5;
                end
              end else if (_T_3291) begin
                release_state <= 3'h1;
              end
            end else if (s2_probe) begin
              if (s2_prb_ack_data) begin
                release_state <= 3'h2;
              end else if (_T_3304) begin
                if (releaseDone) begin
                  release_state <= 3'h7;
                end else begin
                  release_state <= 3'h3;
                end
              end else if (releaseDone) begin
                release_state <= 3'h0;
              end else begin
                release_state <= 3'h5;
              end
            end else if (_T_3291) begin
              release_state <= 3'h1;
            end
          end else if (_T_3308) begin
            if (metaArb_io_in_6_ready) begin
              release_state <= 3'h0;
            end else if (s2_probe) begin
              if (s2_prb_ack_data) begin
                release_state <= 3'h2;
              end else if (_T_3304) begin
                if (releaseDone) begin
                  release_state <= 3'h7;
                end else begin
                  release_state <= 3'h3;
                end
              end else if (releaseDone) begin
                release_state <= 3'h0;
              end else begin
                release_state <= 3'h5;
              end
            end else if (_T_3291) begin
              release_state <= 3'h1;
            end
          end else if (s2_probe) begin
            if (s2_prb_ack_data) begin
              release_state <= 3'h2;
            end else if (_T_3304) begin
              if (releaseDone) begin
                release_state <= 3'h7;
              end else begin
                release_state <= 3'h3;
              end
            end else if (releaseDone) begin
              release_state <= 3'h0;
            end else begin
              release_state <= 3'h5;
            end
          end else if (_T_3291) begin
            release_state <= 3'h1;
          end
        end else if (_T_3312) begin
          if (releaseDone) begin
            release_state <= 3'h0;
          end else if (_T_3308) begin
            if (metaArb_io_in_6_ready) begin
              release_state <= 3'h0;
            end else begin
              release_state <= _GEN_220;
            end
          end else begin
            release_state <= _GEN_220;
          end
        end else if (_T_3308) begin
          if (metaArb_io_in_6_ready) begin
            release_state <= 3'h0;
          end else begin
            release_state <= _GEN_220;
          end
        end else begin
          release_state <= _GEN_220;
        end
      end else if (_T_3313) begin
        if (releaseDone) begin
          release_state <= 3'h7;
        end else if (_T_3312) begin
          if (releaseDone) begin
            release_state <= 3'h0;
          end else begin
            release_state <= _GEN_235;
          end
        end else begin
          release_state <= _GEN_235;
        end
      end else if (_T_3312) begin
        if (releaseDone) begin
          release_state <= 3'h0;
        end else begin
          release_state <= _GEN_235;
        end
      end else begin
        release_state <= _GEN_235;
      end
    end else if (_T_3314) begin
      if (releaseDone) begin
        release_state <= 3'h7;
      end else if (_T_3313) begin
        if (releaseDone) begin
          release_state <= 3'h7;
        end else begin
          release_state <= _GEN_239;
        end
      end else begin
        release_state <= _GEN_239;
      end
    end else if (_T_3313) begin
      if (releaseDone) begin
        release_state <= 3'h7;
      end else begin
        release_state <= _GEN_239;
      end
    end else begin
      release_state <= _GEN_239;
    end
    if (metaReset) begin
      grantInProgress <= 1'h0;
    end else if (reset) begin
      grantInProgress <= 1'h0;
    end else if (_T_3094) begin
      if (grantIsCached) begin
        if (d_last) begin
          grantInProgress <= 1'h0;
        end else begin
          grantInProgress <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      blockProbeAfterGrantCount <= 3'h0;
    end else if (reset) begin
      blockProbeAfterGrantCount <= 3'h0;
    end else if (_T_3094) begin
      if (grantIsCached) begin
        if (d_last) begin
          blockProbeAfterGrantCount <= 3'h7;
        end else if (_T_3224) begin
          blockProbeAfterGrantCount <= _T_3089;
        end
      end else if (_T_3224) begin
        blockProbeAfterGrantCount <= _T_3089;
      end
    end else if (_T_3224) begin
      blockProbeAfterGrantCount <= _T_3089;
    end
    if (metaReset) begin
      lrscCount <= 7'h0;
    end else if (reset) begin
      lrscCount <= 7'h0;
    end else if (s1_probe) begin
      lrscCount <= 7'h0;
    end else if (_T_1269) begin
      lrscCount <= 7'h3;
    end else if (_T_1251) begin
      lrscCount <= _T_1268;
    end else if (_T_1260) begin
      if (s2_hit) begin
        lrscCount <= 7'h4f;
      end else begin
        lrscCount <= 7'h0;
      end
    end
    if (metaReset) begin
      s2_valid_pre_xcpt <= 1'h0;
    end else if (reset) begin
      s2_valid_pre_xcpt <= 1'h0;
    end else begin
      s2_valid_pre_xcpt <= _T_724;
    end
    if (metaReset) begin
      probe_bits_param <= 2'h0;
    end else if (_T_3291) begin
      probe_bits_param <= 2'h0;
    end else if (_T_290) begin
      probe_bits_param <= auto_out_b_bits_param;
    end
    if (metaReset) begin
      probe_bits_size <= 4'h0;
    end else if (_T_3291) begin
      probe_bits_size <= 4'h0;
    end else if (_T_290) begin
      probe_bits_size <= auto_out_b_bits_size;
    end
    if (metaReset) begin
      probe_bits_source <= 1'h0;
    end else if (_T_3291) begin
      probe_bits_source <= 1'h0;
    end else if (_T_290) begin
      probe_bits_source <= auto_out_b_bits_source;
    end
    if (metaReset) begin
      probe_bits_address <= 32'h0;
    end else if (_T_3291) begin
      probe_bits_address <= res_2_address;
    end else if (_T_290) begin
      probe_bits_address <= auto_out_b_bits_address;
    end
    if (metaReset) begin
      s2_probe_state_state <= 2'h0;
    end else if (s1_probe) begin
      s2_probe_state_state <= s1_meta_hit_state_state;
    end
    if (metaReset) begin
      _T_3247 <= 9'h0;
    end else if (reset) begin
      _T_3247 <= 9'h0;
    end else if (_T_3238) begin
      if (c_first) begin
        if (tl_out__c_bits_opcode[0]) begin
          _T_3247 <= _T_3243;
        end else begin
          _T_3247 <= 9'h0;
        end
      end else begin
        _T_3247 <= _T_3250;
      end
    end
    if (metaReset) begin
      s2_release_data_valid <= 1'h0;
    end else begin
      s2_release_data_valid <= s1_release_data_valid & ~releaseRejected;
    end
    if (metaReset) begin
      s1_req_cmd <= 5'h0;
    end else if (s0_clk_en) begin
      s1_req_cmd <= io_cpu_req_bits_cmd;
    end
    if (metaReset) begin
      _T_738 <= 1'h0;
    end else begin
      _T_738 <= ~s1_nack;
    end
    if (metaReset) begin
      s2_req_cmd <= 5'h0;
    end else if (_T_3094) begin
      if (grantIsCached) begin
        if (_T_742) begin
          s2_req_cmd <= s1_req_cmd;
        end
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_cmd <= 5'h0;
        end else if (_T_742) begin
          s2_req_cmd <= s1_req_cmd;
        end
      end else if (_T_742) begin
        s2_req_cmd <= s1_req_cmd;
      end
    end else if (_T_742) begin
      s2_req_cmd <= s1_req_cmd;
    end
    if (metaReset) begin
      s2_hit_state_state <= 2'h0;
    end else if (_T_742) begin
      s2_hit_state_state <= s1_meta_hit_state_state;
    end
    if (metaReset) begin
      lrscAddr <= 34'h0;
    end else if (_T_1260) begin
      lrscAddr <= s2_req_addr[39:6];
    end
    if (metaReset) begin
      s2_req_addr <= 40'h0;
    end else if (_T_3094) begin
      if (grantIsCached) begin
        if (_T_742) begin
          s2_req_addr <= {{8'd0}, tlb_io_resp_paddr};
        end
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_addr <= {{8'd0}, _T_3110};
        end else if (_T_742) begin
          s2_req_addr <= {{8'd0}, tlb_io_resp_paddr};
        end
      end else if (_T_742) begin
        s2_req_addr <= {{8'd0}, tlb_io_resp_paddr};
      end
    end else if (_T_742) begin
      s2_req_addr <= {{8'd0}, tlb_io_resp_paddr};
    end
    if (metaReset) begin
      pstore1_held <= 1'h0;
    end else begin
      pstore1_held <= _T_1470 & ~pstore_drain;
    end
    if (metaReset) begin
      pstore1_addr <= 40'h0;
    end else if (_T_1278) begin
      pstore1_addr <= s1_req_addr;
    end
    if (metaReset) begin
      s1_req_addr <= 40'h0;
    end else if (s0_clk_en) begin
      s1_req_addr <= _T_300;
    end
    if (metaReset) begin
      pstore1_mask <= 8'h0;
    end else if (_T_1278) begin
      if (_T_325) begin
        pstore1_mask <= 8'h0;
      end else begin
        pstore1_mask <= _T_722;
      end
    end
    if (metaReset) begin
      s1_req_typ <= 3'h0;
    end else if (s0_clk_en) begin
      s1_req_typ <= io_cpu_req_bits_typ;
    end
    if (metaReset) begin
      pstore2_valid <= 1'h0;
    end else begin
      pstore2_valid <= _T_1476 | advance_pstore1;
    end
    if (metaReset) begin
      pstore2_addr <= 40'h0;
    end else if (advance_pstore1) begin
      pstore2_addr <= pstore1_addr;
    end
    if (metaReset) begin
      mask <= 8'h0;
    end else if (advance_pstore1) begin
      mask <= pstore1_mask[7:0];
    end
    if (metaReset) begin
      s1_req_tag <= 7'h0;
    end else if (s0_clk_en) begin
      s1_req_tag <= io_cpu_req_bits_tag;
    end
    if (metaReset) begin
      s1_req_phys <= 1'h0;
    end else if (s0_clk_en) begin
      s1_req_phys <= _GEN_9;
    end
    if (metaReset) begin
      s1_flush_valid <= 1'h0;
    end else begin
      s1_flush_valid <= _T_3500 & can_acquire_before_release;
    end
    if (metaReset) begin
      cached_grant_wait <= 1'h0;
    end else if (reset) begin
      cached_grant_wait <= 1'h0;
    end else if (_T_3094) begin
      if (grantIsCached) begin
        if (d_last) begin
          cached_grant_wait <= 1'h0;
        end else if (_T_3058) begin
          if (!(s2_uncached)) begin
            cached_grant_wait <= 1'h1;
          end
        end
      end else if (_T_3058) begin
        if (!(s2_uncached)) begin
          cached_grant_wait <= 1'h1;
        end
      end
    end else if (_T_3058) begin
      if (!(s2_uncached)) begin
        cached_grant_wait <= 1'h1;
      end
    end
    if (metaReset) begin
      release_ack_wait <= 1'h0;
    end else if (reset) begin
      release_ack_wait <= 1'h0;
    end else if (_T_3317) begin
      release_ack_wait <= _GEN_260;
    end else if (_T_3094) begin
      if (!(grantIsCached)) begin
        if (!(grantIsUncached)) begin
          if (grantIsVoluntary) begin
            release_ack_wait <= 1'h0;
          end
        end
      end
    end
    if (metaReset) begin
      uncachedInFlight_0 <= 1'h0;
    end else if (reset) begin
      uncachedInFlight_0 <= 1'h0;
    end else if (_T_3094) begin
      if (grantIsCached) begin
        if (_T_3058) begin
          if (s2_uncached) begin
            uncachedInFlight_0 <= _GEN_99;
          end
        end
      end else if (grantIsUncached) begin
        if (_T_3103) begin
          uncachedInFlight_0 <= 1'h0;
        end else if (_T_3058) begin
          if (s2_uncached) begin
            uncachedInFlight_0 <= _GEN_99;
          end
        end
      end else if (_T_3058) begin
        if (s2_uncached) begin
          uncachedInFlight_0 <= _GEN_99;
        end
      end
    end else if (_T_3058) begin
      if (s2_uncached) begin
        uncachedInFlight_0 <= _GEN_99;
      end
    end
    if (metaReset) begin
      uncachedReqs_0_addr <= 40'h0;
    end else if (_T_3058) begin
      if (s2_uncached) begin
        if (a_sel) begin
          uncachedReqs_0_addr <= s2_req_addr;
        end
      end
    end
    if (metaReset) begin
      uncachedReqs_0_tag <= 7'h0;
    end else if (_T_3058) begin
      if (s2_uncached) begin
        if (a_sel) begin
          uncachedReqs_0_tag <= s2_req_tag;
        end
      end
    end
    if (metaReset) begin
      uncachedReqs_0_typ <= 3'h0;
    end else if (_T_3058) begin
      if (s2_uncached) begin
        if (a_sel) begin
          uncachedReqs_0_typ <= s2_req_typ;
        end
      end
    end
    if (metaReset) begin
      s2_hit_way <= 4'h0;
    end else if (s1_valid_not_nacked) begin
      s2_hit_way <= s1_meta_hit_way;
    end
    if (metaReset) begin
      _T_1060 <= 2'h0;
    end else if (_T_742) begin
      _T_1060 <= s1_victim_way;
    end
    if (metaReset) begin
      s2_probe_way <= 4'h0;
    end else if (s1_probe) begin
      s2_probe_way <= s1_meta_hit_way;
    end
    if (metaReset) begin
      s2_req_tag <= 7'h0;
    end else if (_T_3094) begin
      if (grantIsCached) begin
        if (_T_742) begin
          s2_req_tag <= s1_req_tag;
        end
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_tag <= uncachedReqs_0_tag;
        end else if (_T_742) begin
          s2_req_tag <= s1_req_tag;
        end
      end else if (_T_742) begin
        s2_req_tag <= s1_req_tag;
      end
    end else if (_T_742) begin
      s2_req_tag <= s1_req_tag;
    end
    if (metaReset) begin
      s2_req_typ <= 3'h0;
    end else if (_T_3094) begin
      if (grantIsCached) begin
        if (_T_742) begin
          s2_req_typ <= s1_req_typ;
        end
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_typ <= uncachedReqs_0_typ;
        end else if (_T_742) begin
          s2_req_typ <= s1_req_typ;
        end
      end else if (_T_742) begin
        s2_req_typ <= s1_req_typ;
      end
    end else if (_T_742) begin
      s2_req_typ <= s1_req_typ;
    end
    if (metaReset) begin
      s2_uncached <= 1'h0;
    end else if (_T_742) begin
      s2_uncached <= ~tlb_io_resp_cacheable;
    end
    if (metaReset) begin
      _T_746 <= 40'h0;
    end else if (_T_742) begin
      _T_746 <= s1_req_addr;
    end
    if (metaReset) begin
      s2_flush_valid_pre_tag_ecc <= 1'h0;
    end else begin
      s2_flush_valid_pre_tag_ecc <= s1_flush_valid;
    end
    if (metaReset) begin
      s2_data <= 64'h0;
    end else if (_T_871) begin
      s2_data <= _T_867;
    end
    if (metaReset) begin
      s2_victim_tag <= 20'h0;
    end else if (_T_742) begin
      if (_T_669) begin
        s2_victim_tag <= _T_621[19:0];
      end else if (_T_667) begin
        s2_victim_tag <= _T_614[19:0];
      end else if (_T_665) begin
        s2_victim_tag <= _T_607[19:0];
      end else begin
        s2_victim_tag <= _T_600[19:0];
      end
    end
    if (metaReset) begin
      _T_1068_state <= 2'h0;
    end else if (_T_742) begin
      if (_T_669) begin
        _T_1068_state <= _T_621[21:20];
      end else if (_T_667) begin
        _T_1068_state <= _T_614[21:20];
      end else if (_T_665) begin
        _T_1068_state <= _T_607[21:20];
      end else begin
        _T_1068_state <= _T_600[21:20];
      end
    end
    if (metaReset) begin
      pstore1_cmd <= 5'h0;
    end else if (_T_1278) begin
      pstore1_cmd <= s1_req_cmd;
    end
    if (metaReset) begin
      pstore1_data <= 64'h0;
    end else if (_T_1278) begin
      pstore1_data <= io_cpu_s1_data_data;
    end
    if (metaReset) begin
      pstore1_way <= 4'h0;
    end else if (_T_1278) begin
      pstore1_way <= s1_meta_hit_way;
    end
    if (metaReset) begin
      pstore1_rmw <= 1'h0;
    end else if (_T_1278) begin
      pstore1_rmw <= _T_1340;
    end
    if (metaReset) begin
      pstore2_way <= 4'h0;
    end else if (advance_pstore1) begin
      pstore2_way <= pstore1_way;
    end
    if (metaReset) begin
      _T_1487 <= 8'h0;
    end else if (advance_pstore1) begin
      _T_1487 <= pstore1_storegen_data[7:0];
    end
    if (metaReset) begin
      _T_1493 <= 8'h0;
    end else if (advance_pstore1) begin
      _T_1493 <= pstore1_storegen_data[15:8];
    end
    if (metaReset) begin
      _T_1499 <= 8'h0;
    end else if (advance_pstore1) begin
      _T_1499 <= pstore1_storegen_data[23:16];
    end
    if (metaReset) begin
      _T_1505 <= 8'h0;
    end else if (advance_pstore1) begin
      _T_1505 <= pstore1_storegen_data[31:24];
    end
    if (metaReset) begin
      _T_1511 <= 8'h0;
    end else if (advance_pstore1) begin
      _T_1511 <= pstore1_storegen_data[39:32];
    end
    if (metaReset) begin
      _T_1517 <= 8'h0;
    end else if (advance_pstore1) begin
      _T_1517 <= pstore1_storegen_data[47:40];
    end
    if (metaReset) begin
      _T_1523 <= 8'h0;
    end else if (advance_pstore1) begin
      _T_1523 <= pstore1_storegen_data[55:48];
    end
    if (metaReset) begin
      _T_1529 <= 8'h0;
    end else if (advance_pstore1) begin
      _T_1529 <= pstore1_storegen_data[63:56];
    end
    if (metaReset) begin
      s1_release_data_valid <= 1'h0;
    end else begin
      s1_release_data_valid <= dataArb_io_in_2_ready & dataArb_io_in_2_valid;
    end
    if (metaReset) begin
      _T_3374 <= 1'h0;
    end else begin
      _T_3374 <= tlb_io_req_valid & ~s1_nack;
    end
    if (metaReset) begin
      _T_3376_pf_ld <= 1'h0;
    end else if (s1_valid_not_nacked) begin
      _T_3376_pf_ld <= tlb_io_resp_pf_ld;
    end
    if (metaReset) begin
      _T_3376_pf_st <= 1'h0;
    end else if (s1_valid_not_nacked) begin
      _T_3376_pf_st <= tlb_io_resp_pf_st;
    end
    if (metaReset) begin
      _T_3376_ae_ld <= 1'h0;
    end else if (s1_valid_not_nacked) begin
      _T_3376_ae_ld <= tlb_io_resp_ae_ld;
    end
    if (metaReset) begin
      _T_3376_ae_st <= 1'h0;
    end else if (s1_valid_not_nacked) begin
      _T_3376_ae_st <= tlb_io_resp_ae_st;
    end
    if (metaReset) begin
      _T_3376_ma_ld <= 1'h0;
    end else if (s1_valid_not_nacked) begin
      _T_3376_ma_ld <= tlb_io_resp_ma_ld;
    end
    if (metaReset) begin
      _T_3376_ma_st <= 1'h0;
    end else if (s1_valid_not_nacked) begin
      _T_3376_ma_st <= tlb_io_resp_ma_st;
    end
    if (metaReset) begin
      doUncachedResp <= 1'h0;
    end else begin
      doUncachedResp <= io_cpu_replay_next;
    end
    if (metaReset) begin
      resetting <= 1'h0;
    end else if (reset) begin
      resetting <= 1'h0;
    end else if (resetting) begin
      if (flushDone) begin
        resetting <= 1'h0;
      end else begin
        resetting <= _GEN_290;
      end
    end else begin
      resetting <= _GEN_290;
    end
    if (metaReset) begin
      _T_3473 <= 1'h0;
    end else begin
      _T_3473 <= reset;
    end
    if (metaReset) begin
      flushed <= 1'h0;
    end else begin
      flushed <= reset | flushed;
    end
    if (metaReset) begin
      flushing <= 1'h0;
    end else if (reset) begin
      flushing <= 1'h0;
    end else if (_T_3479) begin
      if (~flushed) begin
        flushing <= _T_3487;
      end
    end
    if (metaReset) begin
      flushCounter <= 8'h0;
    end else if (reset) begin
      flushCounter <= 8'hc0;
    end else begin
      flushCounter <= _GEN_295[7:0];
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_471) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:913 assert(!needsRead(req) || res)\n"); // @[DCache.scala 913:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_471) begin
          $fatal; // @[DCache.scala 913:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_471) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:913 assert(!needsRead(req) || res)\n"); // @[DCache.scala 913:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_471) begin
          $fatal; // @[DCache.scala 913:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_1441) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:366 assert(pstore1_rmw || pstore1_valid_not_rmw(io.cpu.s2_kill) === pstore1_valid)\n"); // @[DCache.scala 366:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_1441) begin
          $fatal; // @[DCache.scala 366:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_308 & ~_T_3096) begin
          $fwrite(32'h80000002,"Assertion failed: A GrantData was unexpected by the dcache.\n    at DCache.scala:500 assert(cached_grant_wait, \"A GrantData was unexpected by the dcache.\")\n"); // @[DCache.scala 500:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_308 & ~_T_3096) begin
          $fatal; // @[DCache.scala 500:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_313 & ~_T_3105) begin
          $fwrite(32'h80000002,"Assertion failed: An AccessAck was unexpected by the dcache.\n    at DCache.scala:512 assert(f, \"An AccessAck was unexpected by the dcache.\") // TODO must handle Ack coming back on same cycle!\n"); // @[DCache.scala 512:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_313 & ~_T_3105) begin
          $fatal; // @[DCache.scala 512:17]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_322 & ~_T_3112) begin
          $fwrite(32'h80000002,"Assertion failed: A ReleaseAck was unexpected by the dcache.\n    at DCache.scala:530 assert(release_ack_wait, \"A ReleaseAck was unexpected by the dcache.\") // TODO should handle Ack coming back on same cycle!\n"); // @[DCache.scala 530:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_322 & ~_T_3112) begin
          $fatal; // @[DCache.scala 530:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_3125) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:538 assert(tl_out.e.fire() === (tl_out.d.fire() && d_first && grantIsCached))\n"); // @[DCache.scala 538:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_3125) begin
          $fatal; // @[DCache.scala 538:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3291 & ~_T_3297) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:616 assert(!(s2_valid && s2_hit_valid && !s2_data_error))\n"); // @[DCache.scala 616:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3291 & ~_T_3297) begin
          $fatal; // @[DCache.scala 616:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (doUncachedResp & ~_T_3403) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:723 assert(!s2_valid_hit)\n"); // @[DCache.scala 723:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (doUncachedResp & ~_T_3403) begin
          $fatal; // @[DCache.scala 723:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    DCache_state <= DCache_xor0;
    if (!(DCache_cov_read_data)) begin
      DCache_covSum <= DCache_covSum + 1'h1;
    end
  end
  always @(posedge gated_clock) begin
    if(DCache_cov_write_en & DCache_cov_write_mask) begin
      DCache_cov[DCache_cov_write_addr] <= DCache_cov_write_data; // @[Coverage map for DCache]
    end
  end
endmodule
module Frontend(
  input         gated_clock,
  input         reset,
  input         auto_icache_master_out_a_ready,
  output        auto_icache_master_out_a_valid,
  output [31:0] auto_icache_master_out_a_bits_address,
  input         auto_icache_master_out_d_valid,
  input  [2:0]  auto_icache_master_out_d_bits_opcode,
  input  [3:0]  auto_icache_master_out_d_bits_size,
  input  [63:0] auto_icache_master_out_d_bits_data,
  input         auto_icache_master_out_d_bits_corrupt,
  input  [31:0] io_reset_vector,
  input         io_cpu_might_request,
  input         io_cpu_req_valid,
  input  [39:0] io_cpu_req_bits_pc,
  input         io_cpu_req_bits_speculative,
  input         io_cpu_sfence_valid,
  input         io_cpu_sfence_bits_rs1,
  input         io_cpu_sfence_bits_rs2,
  input  [38:0] io_cpu_sfence_bits_addr,
  input         io_cpu_resp_ready,
  output        io_cpu_resp_valid,
  output        io_cpu_resp_bits_btb_taken,
  output        io_cpu_resp_bits_btb_bridx,
  output [4:0]  io_cpu_resp_bits_btb_entry,
  output [7:0]  io_cpu_resp_bits_btb_bht_history,
  output [39:0] io_cpu_resp_bits_pc,
  output [31:0] io_cpu_resp_bits_data,
  output        io_cpu_resp_bits_xcpt_pf_inst,
  output        io_cpu_resp_bits_xcpt_ae_inst,
  output        io_cpu_resp_bits_replay,
  input         io_cpu_btb_update_valid,
  input  [4:0]  io_cpu_btb_update_bits_prediction_entry,
  input  [38:0] io_cpu_btb_update_bits_pc,
  input         io_cpu_btb_update_bits_isValid,
  input  [38:0] io_cpu_btb_update_bits_br_pc,
  input  [1:0]  io_cpu_btb_update_bits_cfiType,
  input         io_cpu_bht_update_valid,
  input  [7:0]  io_cpu_bht_update_bits_prediction_history,
  input  [38:0] io_cpu_bht_update_bits_pc,
  input         io_cpu_bht_update_bits_branch,
  input         io_cpu_bht_update_bits_taken,
  input         io_cpu_bht_update_bits_mispredict,
  input         io_cpu_flush_icache,
  output [39:0] io_cpu_npc,
  input         io_ptw_req_ready,
  output        io_ptw_req_valid,
  output        io_ptw_req_bits_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  input         io_ptw_resp_valid,
  input         io_ptw_resp_bits_ae,
  input  [53:0] io_ptw_resp_bits_pte_ppn,
  input         io_ptw_resp_bits_pte_d,
  input         io_ptw_resp_bits_pte_a,
  input         io_ptw_resp_bits_pte_g,
  input         io_ptw_resp_bits_pte_u,
  input         io_ptw_resp_bits_pte_x,
  input         io_ptw_resp_bits_pte_w,
  input         io_ptw_resp_bits_pte_r,
  input         io_ptw_resp_bits_pte_v,
  input  [1:0]  io_ptw_resp_bits_level,
  input         io_ptw_resp_bits_homogeneous,
  input  [3:0]  io_ptw_ptbr_mode,
  input  [1:0]  io_ptw_status_prv,
  input         io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
  input         io_ptw_pmp_0_cfg_w,
  input         io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr,
  input  [31:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
  input         io_ptw_pmp_1_cfg_w,
  input         io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr,
  input  [31:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
  input         io_ptw_pmp_2_cfg_w,
  input         io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr,
  input  [31:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
  input         io_ptw_pmp_3_cfg_w,
  input         io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr,
  input  [31:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
  input         io_ptw_pmp_4_cfg_w,
  input         io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr,
  input  [31:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
  input         io_ptw_pmp_5_cfg_w,
  input         io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr,
  input  [31:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
  input         io_ptw_pmp_6_cfg_w,
  input         io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr,
  input  [31:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
  input         io_ptw_pmp_7_cfg_w,
  input         io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr,
  input  [31:0] io_ptw_pmp_7_mask,
  input  [26:0] io_ptw_vpoffset_bits_value,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         icache_halt,
  input         fq_halt,
  input         tlb_halt,
  input         btb_halt
);
  wire  icache_clock; // @[Frontend.scala 61:26]
  wire  icache_reset; // @[Frontend.scala 61:26]
  wire  icache_auto_master_out_a_ready; // @[Frontend.scala 61:26]
  wire  icache_auto_master_out_a_valid; // @[Frontend.scala 61:26]
  wire [31:0] icache_auto_master_out_a_bits_address; // @[Frontend.scala 61:26]
  wire  icache_auto_master_out_d_valid; // @[Frontend.scala 61:26]
  wire [2:0] icache_auto_master_out_d_bits_opcode; // @[Frontend.scala 61:26]
  wire [3:0] icache_auto_master_out_d_bits_size; // @[Frontend.scala 61:26]
  wire [63:0] icache_auto_master_out_d_bits_data; // @[Frontend.scala 61:26]
  wire  icache_auto_master_out_d_bits_corrupt; // @[Frontend.scala 61:26]
  wire  icache_io_req_ready; // @[Frontend.scala 61:26]
  wire  icache_io_req_valid; // @[Frontend.scala 61:26]
  wire [38:0] icache_io_req_bits_addr; // @[Frontend.scala 61:26]
  wire [31:0] icache_io_s1_paddr; // @[Frontend.scala 61:26]
  wire  icache_io_s1_kill; // @[Frontend.scala 61:26]
  wire  icache_io_s2_kill; // @[Frontend.scala 61:26]
  wire  icache_io_resp_valid; // @[Frontend.scala 61:26]
  wire [31:0] icache_io_resp_bits_data; // @[Frontend.scala 61:26]
  wire  icache_io_resp_bits_ae; // @[Frontend.scala 61:26]
  wire  icache_io_invalidate; // @[Frontend.scala 61:26]
  wire [29:0] icache_io_covSum; // @[Frontend.scala 61:26]
  wire  icache_metaAssert; // @[Frontend.scala 61:26]
  wire  icache_metaReset; // @[Frontend.scala 61:26]
  wire  fq_clock; // @[Frontend.scala 82:57]
  wire  fq_reset; // @[Frontend.scala 82:57]
  wire  fq_io_enq_ready; // @[Frontend.scala 82:57]
  wire  fq_io_enq_valid; // @[Frontend.scala 82:57]
  wire  fq_io_enq_bits_btb_taken; // @[Frontend.scala 82:57]
  wire  fq_io_enq_bits_btb_bridx; // @[Frontend.scala 82:57]
  wire [4:0] fq_io_enq_bits_btb_entry; // @[Frontend.scala 82:57]
  wire [7:0] fq_io_enq_bits_btb_bht_history; // @[Frontend.scala 82:57]
  wire [39:0] fq_io_enq_bits_pc; // @[Frontend.scala 82:57]
  wire [31:0] fq_io_enq_bits_data; // @[Frontend.scala 82:57]
  wire [1:0] fq_io_enq_bits_mask; // @[Frontend.scala 82:57]
  wire  fq_io_enq_bits_xcpt_pf_inst; // @[Frontend.scala 82:57]
  wire  fq_io_enq_bits_xcpt_ae_inst; // @[Frontend.scala 82:57]
  wire  fq_io_enq_bits_replay; // @[Frontend.scala 82:57]
  wire  fq_io_deq_ready; // @[Frontend.scala 82:57]
  wire  fq_io_deq_valid; // @[Frontend.scala 82:57]
  wire  fq_io_deq_bits_btb_taken; // @[Frontend.scala 82:57]
  wire  fq_io_deq_bits_btb_bridx; // @[Frontend.scala 82:57]
  wire [4:0] fq_io_deq_bits_btb_entry; // @[Frontend.scala 82:57]
  wire [7:0] fq_io_deq_bits_btb_bht_history; // @[Frontend.scala 82:57]
  wire [39:0] fq_io_deq_bits_pc; // @[Frontend.scala 82:57]
  wire [31:0] fq_io_deq_bits_data; // @[Frontend.scala 82:57]
  wire  fq_io_deq_bits_xcpt_pf_inst; // @[Frontend.scala 82:57]
  wire  fq_io_deq_bits_xcpt_ae_inst; // @[Frontend.scala 82:57]
  wire  fq_io_deq_bits_replay; // @[Frontend.scala 82:57]
  wire [4:0] fq_io_mask; // @[Frontend.scala 82:57]
  wire [29:0] fq_io_covSum; // @[Frontend.scala 82:57]
  wire  fq_metaAssert; // @[Frontend.scala 82:57]
  wire  fq_metaReset; // @[Frontend.scala 82:57]
  wire  tlb_clock; // @[Frontend.scala 95:19]
  wire  tlb_reset; // @[Frontend.scala 95:19]
  wire  tlb_io_req_ready; // @[Frontend.scala 95:19]
  wire  tlb_io_req_valid; // @[Frontend.scala 95:19]
  wire [39:0] tlb_io_req_bits_vaddr; // @[Frontend.scala 95:19]
  wire  tlb_io_resp_miss; // @[Frontend.scala 95:19]
  wire [31:0] tlb_io_resp_paddr; // @[Frontend.scala 95:19]
  wire  tlb_io_resp_pf_inst; // @[Frontend.scala 95:19]
  wire  tlb_io_resp_ae_inst; // @[Frontend.scala 95:19]
  wire  tlb_io_resp_cacheable; // @[Frontend.scala 95:19]
  wire  tlb_io_sfence_valid; // @[Frontend.scala 95:19]
  wire  tlb_io_sfence_bits_rs1; // @[Frontend.scala 95:19]
  wire  tlb_io_sfence_bits_rs2; // @[Frontend.scala 95:19]
  wire [38:0] tlb_io_sfence_bits_addr; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_req_ready; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_req_valid; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_req_bits_valid; // @[Frontend.scala 95:19]
  wire [26:0] tlb_io_ptw_req_bits_bits_addr; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_resp_valid; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_resp_bits_ae; // @[Frontend.scala 95:19]
  wire [53:0] tlb_io_ptw_resp_bits_pte_ppn; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_resp_bits_pte_d; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_resp_bits_pte_a; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_resp_bits_pte_g; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_resp_bits_pte_u; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_resp_bits_pte_x; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_resp_bits_pte_w; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_resp_bits_pte_r; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_resp_bits_pte_v; // @[Frontend.scala 95:19]
  wire [1:0] tlb_io_ptw_resp_bits_level; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_resp_bits_homogeneous; // @[Frontend.scala 95:19]
  wire [3:0] tlb_io_ptw_ptbr_mode; // @[Frontend.scala 95:19]
  wire [1:0] tlb_io_ptw_status_prv; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_0_cfg_l; // @[Frontend.scala 95:19]
  wire [1:0] tlb_io_ptw_pmp_0_cfg_a; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_0_cfg_x; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_0_cfg_w; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_0_cfg_r; // @[Frontend.scala 95:19]
  wire [29:0] tlb_io_ptw_pmp_0_addr; // @[Frontend.scala 95:19]
  wire [31:0] tlb_io_ptw_pmp_0_mask; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_1_cfg_l; // @[Frontend.scala 95:19]
  wire [1:0] tlb_io_ptw_pmp_1_cfg_a; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_1_cfg_x; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_1_cfg_w; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_1_cfg_r; // @[Frontend.scala 95:19]
  wire [29:0] tlb_io_ptw_pmp_1_addr; // @[Frontend.scala 95:19]
  wire [31:0] tlb_io_ptw_pmp_1_mask; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_2_cfg_l; // @[Frontend.scala 95:19]
  wire [1:0] tlb_io_ptw_pmp_2_cfg_a; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_2_cfg_x; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_2_cfg_w; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_2_cfg_r; // @[Frontend.scala 95:19]
  wire [29:0] tlb_io_ptw_pmp_2_addr; // @[Frontend.scala 95:19]
  wire [31:0] tlb_io_ptw_pmp_2_mask; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_3_cfg_l; // @[Frontend.scala 95:19]
  wire [1:0] tlb_io_ptw_pmp_3_cfg_a; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_3_cfg_x; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_3_cfg_w; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_3_cfg_r; // @[Frontend.scala 95:19]
  wire [29:0] tlb_io_ptw_pmp_3_addr; // @[Frontend.scala 95:19]
  wire [31:0] tlb_io_ptw_pmp_3_mask; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_4_cfg_l; // @[Frontend.scala 95:19]
  wire [1:0] tlb_io_ptw_pmp_4_cfg_a; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_4_cfg_x; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_4_cfg_w; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_4_cfg_r; // @[Frontend.scala 95:19]
  wire [29:0] tlb_io_ptw_pmp_4_addr; // @[Frontend.scala 95:19]
  wire [31:0] tlb_io_ptw_pmp_4_mask; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_5_cfg_l; // @[Frontend.scala 95:19]
  wire [1:0] tlb_io_ptw_pmp_5_cfg_a; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_5_cfg_x; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_5_cfg_w; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_5_cfg_r; // @[Frontend.scala 95:19]
  wire [29:0] tlb_io_ptw_pmp_5_addr; // @[Frontend.scala 95:19]
  wire [31:0] tlb_io_ptw_pmp_5_mask; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_6_cfg_l; // @[Frontend.scala 95:19]
  wire [1:0] tlb_io_ptw_pmp_6_cfg_a; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_6_cfg_x; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_6_cfg_w; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_6_cfg_r; // @[Frontend.scala 95:19]
  wire [29:0] tlb_io_ptw_pmp_6_addr; // @[Frontend.scala 95:19]
  wire [31:0] tlb_io_ptw_pmp_6_mask; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_7_cfg_l; // @[Frontend.scala 95:19]
  wire [1:0] tlb_io_ptw_pmp_7_cfg_a; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_7_cfg_x; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_7_cfg_w; // @[Frontend.scala 95:19]
  wire  tlb_io_ptw_pmp_7_cfg_r; // @[Frontend.scala 95:19]
  wire [29:0] tlb_io_ptw_pmp_7_addr; // @[Frontend.scala 95:19]
  wire [31:0] tlb_io_ptw_pmp_7_mask; // @[Frontend.scala 95:19]
  wire [26:0] tlb_io_ptw_vpoffset_bits_value; // @[Frontend.scala 95:19]
  wire  tlb_io_kill; // @[Frontend.scala 95:19]
  wire [29:0] tlb_io_covSum; // @[Frontend.scala 95:19]
  wire  tlb_metaAssert; // @[Frontend.scala 95:19]
  wire  tlb_metaReset; // @[Frontend.scala 95:19]
  wire  btb_clock; // @[Frontend.scala 170:21]
  wire  btb_reset; // @[Frontend.scala 170:21]
  wire [38:0] btb_io_req_bits_addr; // @[Frontend.scala 170:21]
  wire  btb_io_resp_valid; // @[Frontend.scala 170:21]
  wire  btb_io_resp_bits_taken; // @[Frontend.scala 170:21]
  wire  btb_io_resp_bits_bridx; // @[Frontend.scala 170:21]
  wire [38:0] btb_io_resp_bits_target; // @[Frontend.scala 170:21]
  wire [4:0] btb_io_resp_bits_entry; // @[Frontend.scala 170:21]
  wire [7:0] btb_io_resp_bits_bht_history; // @[Frontend.scala 170:21]
  wire  btb_io_resp_bits_bht_value; // @[Frontend.scala 170:21]
  wire  btb_io_btb_update_valid; // @[Frontend.scala 170:21]
  wire [4:0] btb_io_btb_update_bits_prediction_entry; // @[Frontend.scala 170:21]
  wire [38:0] btb_io_btb_update_bits_pc; // @[Frontend.scala 170:21]
  wire  btb_io_btb_update_bits_isValid; // @[Frontend.scala 170:21]
  wire [38:0] btb_io_btb_update_bits_br_pc; // @[Frontend.scala 170:21]
  wire [1:0] btb_io_btb_update_bits_cfiType; // @[Frontend.scala 170:21]
  wire  btb_io_bht_update_valid; // @[Frontend.scala 170:21]
  wire [7:0] btb_io_bht_update_bits_prediction_history; // @[Frontend.scala 170:21]
  wire [38:0] btb_io_bht_update_bits_pc; // @[Frontend.scala 170:21]
  wire  btb_io_bht_update_bits_branch; // @[Frontend.scala 170:21]
  wire  btb_io_bht_update_bits_taken; // @[Frontend.scala 170:21]
  wire  btb_io_bht_update_bits_mispredict; // @[Frontend.scala 170:21]
  wire  btb_io_bht_advance_valid; // @[Frontend.scala 170:21]
  wire  btb_io_bht_advance_bits_bht_value; // @[Frontend.scala 170:21]
  wire  btb_io_ras_update_valid; // @[Frontend.scala 170:21]
  wire [1:0] btb_io_ras_update_bits_cfiType; // @[Frontend.scala 170:21]
  wire [38:0] btb_io_ras_update_bits_returnAddr; // @[Frontend.scala 170:21]
  wire  btb_io_ras_head_valid; // @[Frontend.scala 170:21]
  wire [38:0] btb_io_ras_head_bits; // @[Frontend.scala 170:21]
  wire  btb_io_flush; // @[Frontend.scala 170:21]
  wire [29:0] btb_io_covSum; // @[Frontend.scala 170:21]
  wire  btb_metaAssert; // @[Frontend.scala 170:21]
  wire  btb_metaReset; // @[Frontend.scala 170:21]
  wire  _T_212; // @[Frontend.scala 86:29]
  wire  _T_213; // @[Frontend.scala 86:52]
  wire  _T_214; // @[Frontend.scala 86:75]
  wire  _T_215; // @[Frontend.scala 86:102]
  wire  _T_217; // @[Frontend.scala 86:130]
  wire  _T_219; // @[Frontend.scala 86:9]
  wire  s0_valid; // @[Frontend.scala 97:35]
  reg  s1_valid; // @[Frontend.scala 98:25]
  reg [31:0] _RAND_0;
  reg [39:0] s1_pc; // @[Frontend.scala 99:18]
  reg [63:0] _RAND_1;
  reg  s1_speculative; // @[Frontend.scala 100:27]
  reg [31:0] _RAND_2;
  reg  s2_valid; // @[Frontend.scala 101:25]
  reg [31:0] _RAND_3;
  wire [31:0] _T_229; // @[Frontend.scala 331:33]
  reg [39:0] s2_pc; // @[Frontend.scala 102:22]
  reg [63:0] _RAND_4;
  reg  s2_btb_resp_valid; // @[Frontend.scala 103:44]
  reg [31:0] _RAND_5;
  reg  s2_btb_resp_bits_taken; // @[Frontend.scala 104:29]
  reg [31:0] _RAND_6;
  reg  s2_btb_resp_bits_bridx; // @[Frontend.scala 104:29]
  reg [31:0] _RAND_7;
  reg [4:0] s2_btb_resp_bits_entry; // @[Frontend.scala 104:29]
  reg [31:0] _RAND_8;
  reg [7:0] s2_btb_resp_bits_bht_history; // @[Frontend.scala 104:29]
  reg [31:0] _RAND_9;
  reg  s2_btb_resp_bits_bht_value; // @[Frontend.scala 104:29]
  reg [31:0] _RAND_10;
  wire  s2_btb_taken; // @[Frontend.scala 105:40]
  reg  s2_tlb_resp_miss; // @[Frontend.scala 106:24]
  reg [31:0] _RAND_11;
  reg  s2_tlb_resp_pf_inst; // @[Frontend.scala 106:24]
  reg [31:0] _RAND_12;
  reg  s2_tlb_resp_ae_inst; // @[Frontend.scala 106:24]
  reg [31:0] _RAND_13;
  reg  s2_tlb_resp_cacheable; // @[Frontend.scala 106:24]
  reg [31:0] _RAND_14;
  wire  s2_xcpt; // @[Frontend.scala 107:37]
  reg  s2_speculative; // @[Frontend.scala 108:27]
  reg [31:0] _RAND_15;
  reg  s2_partial_insn_valid; // @[Frontend.scala 109:38]
  reg [31:0] _RAND_16;
  reg [15:0] s2_partial_insn; // @[Frontend.scala 110:28]
  reg [31:0] _RAND_17;
  reg  wrong_path; // @[Frontend.scala 111:23]
  reg [31:0] _RAND_18;
  wire [39:0] _T_238; // @[Frontend.scala 113:29]
  wire [39:0] s1_base_pc; // @[Frontend.scala 113:20]
  wire [39:0] ntpc; // @[Frontend.scala 114:25]
  wire  _T_243; // @[Decoupled.scala 37:37]
  wire  _T_245; // @[Frontend.scala 119:26]
  reg  _T_249; // @[Frontend.scala 119:58]
  reg [31:0] _RAND_19;
  wire  s2_replay; // @[Frontend.scala 119:48]
  wire  _T_247; // @[Frontend.scala 119:69]
  wire  _T_310; // @[Frontend.scala 199:45]
  wire  taken_prevRVI; // @[Frontend.scala 200:31]
  wire [15:0] taken_bits; // @[Frontend.scala 202:37]
  wire [31:0] taken_rviBits; // @[Cat.scala 30:58]
  wire  taken_rviJump; // @[Frontend.scala 206:34]
  wire  taken_rviJALR; // @[Frontend.scala 207:34]
  wire  _T_504; // @[Frontend.scala 221:29]
  wire  taken_rviBranch; // @[Frontend.scala 205:36]
  wire  _T_505; // @[Frontend.scala 221:53]
  wire  _T_506; // @[Frontend.scala 221:40]
  wire  _T_507; // @[Frontend.scala 221:17]
  wire  taken_valid; // @[Frontend.scala 201:44]
  wire [15:0] _T_332; // @[Frontend.scala 212:26]
  wire  taken_rvcJump; // @[Frontend.scala 212:26]
  wire [15:0] _T_374; // @[Frontend.scala 216:26]
  wire  _T_375; // @[Frontend.scala 216:26]
  wire  _T_377; // @[Frontend.scala 216:62]
  wire  taken_rvcJALR; // @[Frontend.scala 216:49]
  wire  _T_508; // @[Frontend.scala 222:27]
  wire  _T_368; // @[Frontend.scala 214:24]
  wire  taken_rvcJR; // @[Frontend.scala 214:46]
  wire  _T_509; // @[Frontend.scala 222:38]
  wire  _T_327; // @[Frontend.scala 210:28]
  wire  _T_329; // @[Frontend.scala 210:60]
  wire  taken_rvcBranch; // @[Frontend.scala 210:52]
  wire  _T_510; // @[Frontend.scala 222:60]
  wire  _T_511; // @[Frontend.scala 222:47]
  wire  _T_512; // @[Frontend.scala 222:15]
  wire  taken_taken; // @[Frontend.scala 221:71]
  wire  taken_idx; // @[Frontend.scala 236:13]
  wire  _T_577; // @[Frontend.scala 199:45]
  wire  taken_prevRVI_1; // @[Frontend.scala 200:31]
  wire [15:0] taken_bits_1; // @[Frontend.scala 202:37]
  wire [31:0] taken_rviBits_1; // @[Cat.scala 30:58]
  wire  taken_rviJALR_1; // @[Frontend.scala 207:34]
  wire  _T_587; // @[Frontend.scala 208:31]
  wire [4:0] _T_589; // @[Frontend.scala 208:66]
  wire  _T_590; // @[Frontend.scala 208:66]
  wire  taken_rviReturn_1; // @[Frontend.scala 208:46]
  wire  _T_780; // @[Frontend.scala 223:61]
  wire  taken_valid_1; // @[Frontend.scala 201:44]
  wire [15:0] _T_634; // @[Frontend.scala 214:24]
  wire  _T_635; // @[Frontend.scala 214:24]
  wire  _T_637; // @[Frontend.scala 214:59]
  wire  taken_rvcJR_1; // @[Frontend.scala 214:46]
  wire [4:0] _T_639; // @[Frontend.scala 215:49]
  wire  _T_640; // @[Frontend.scala 215:49]
  wire  taken_rvcReturn_1; // @[Frontend.scala 215:29]
  wire  _T_781; // @[Frontend.scala 223:83]
  wire  _T_782; // @[Frontend.scala 223:74]
  wire  taken_predictReturn_1; // @[Frontend.scala 223:49]
  wire  _T_821; // @[Frontend.scala 249:26]
  wire  _T_320; // @[Frontend.scala 208:31]
  wire [4:0] _T_322; // @[Frontend.scala 208:66]
  wire  _T_323; // @[Frontend.scala 208:66]
  wire  taken_rviReturn; // @[Frontend.scala 208:46]
  wire  _T_513; // @[Frontend.scala 223:61]
  wire [4:0] _T_372; // @[Frontend.scala 215:49]
  wire  _T_373; // @[Frontend.scala 215:49]
  wire  taken_rvcReturn; // @[Frontend.scala 215:29]
  wire  _T_514; // @[Frontend.scala 223:83]
  wire  _T_515; // @[Frontend.scala 223:74]
  wire  taken_predictReturn; // @[Frontend.scala 223:49]
  wire  _T_554; // @[Frontend.scala 249:26]
  wire  _GEN_44; // @[Frontend.scala 245:30]
  wire  _GEN_77; // @[Frontend.scala 249:44]
  wire  _GEN_80; // @[Frontend.scala 245:30]
  wire  useRAS; // @[Frontend.scala 236:25]
  wire  taken_rviBranch_1; // @[Frontend.scala 205:36]
  wire  _T_785; // @[Frontend.scala 225:53]
  wire [15:0] _T_593; // @[Frontend.scala 210:28]
  wire  _T_594; // @[Frontend.scala 210:28]
  wire  _T_596; // @[Frontend.scala 210:60]
  wire  taken_rvcBranch_1; // @[Frontend.scala 210:52]
  wire  _T_786; // @[Frontend.scala 225:75]
  wire  _T_787; // @[Frontend.scala 225:66]
  wire  taken_predictBranch_1; // @[Frontend.scala 225:41]
  wire  taken_rviJump_1; // @[Frontend.scala 206:34]
  wire  _T_783; // @[Frontend.scala 224:33]
  wire  taken_rvcJump_1; // @[Frontend.scala 212:26]
  wire  _T_784; // @[Frontend.scala 224:53]
  wire  taken_predictJump_1; // @[Frontend.scala 224:44]
  wire  _T_822; // @[Frontend.scala 252:44]
  wire  _T_823; // @[Frontend.scala 252:26]
  wire [39:0] _T_292; // @[Frontend.scala 192:31]
  wire [39:0] s2_base_pc; // @[Frontend.scala 192:22]
  wire [39:0] taken_pc_1; // @[Frontend.scala 253:33]
  wire [39:0] _T_826; // @[Frontend.scala 256:36]
  wire [39:0] _T_828; // @[Frontend.scala 256:57]
  wire  _T_648; // @[RocketCore.scala 954:53]
  wire  _T_703; // @[Cat.scala 30:58]
  wire [10:0] _T_702; // @[Cat.scala 30:58]
  wire [7:0] _T_700; // @[Cat.scala 30:58]
  wire  _T_699; // @[Cat.scala 30:58]
  wire [31:0] _T_707; // @[RocketCore.scala 968:53]
  wire [7:0] _T_762; // @[Cat.scala 30:58]
  wire  _T_761; // @[Cat.scala 30:58]
  wire [31:0] _T_769; // @[RocketCore.scala 968:53]
  wire [31:0] taken_rviImm_1; // @[Frontend.scala 218:23]
  wire [4:0] _T_604; // @[Bitwise.scala 72:12]
  wire [12:0] _T_614; // @[Frontend.scala 213:66]
  wire [9:0] _T_617; // @[Bitwise.scala 72:12]
  wire [20:0] _T_633; // @[Frontend.scala 213:106]
  wire [20:0] taken_rvcImm_1; // @[Frontend.scala 213:23]
  wire [31:0] _T_829; // @[Frontend.scala 256:69]
  wire [39:0] _GEN_126; // @[Frontend.scala 256:64]
  wire [39:0] _T_832; // @[Frontend.scala 257:34]
  wire  _T_518; // @[Frontend.scala 225:53]
  wire  _T_519; // @[Frontend.scala 225:75]
  wire  _T_520; // @[Frontend.scala 225:66]
  wire  taken_predictBranch; // @[Frontend.scala 225:41]
  wire  _T_516; // @[Frontend.scala 224:33]
  wire  _T_517; // @[Frontend.scala 224:53]
  wire  taken_predictJump; // @[Frontend.scala 224:44]
  wire  _T_555; // @[Frontend.scala 252:44]
  wire  _T_556; // @[Frontend.scala 252:26]
  wire [39:0] _T_557; // @[Frontend.scala 255:32]
  wire  _T_381; // @[RocketCore.scala 954:53]
  wire  _T_436; // @[Cat.scala 30:58]
  wire [10:0] _T_435; // @[Cat.scala 30:58]
  wire [7:0] _T_433; // @[Cat.scala 30:58]
  wire  _T_432; // @[Cat.scala 30:58]
  wire [31:0] _T_440; // @[RocketCore.scala 968:53]
  wire [7:0] _T_495; // @[Cat.scala 30:58]
  wire  _T_494; // @[Cat.scala 30:58]
  wire [31:0] _T_502; // @[RocketCore.scala 968:53]
  wire [31:0] taken_rviImm; // @[Frontend.scala 218:23]
  wire [32:0] _T_558; // @[Frontend.scala 255:61]
  wire [4:0] _T_337; // @[Bitwise.scala 72:12]
  wire [12:0] _T_347; // @[Frontend.scala 213:66]
  wire [9:0] _T_350; // @[Bitwise.scala 72:12]
  wire [20:0] _T_366; // @[Frontend.scala 213:106]
  wire [20:0] taken_rvcImm; // @[Frontend.scala 213:23]
  wire [32:0] _T_559; // @[Frontend.scala 255:44]
  wire [39:0] _GEN_127; // @[Frontend.scala 255:39]
  wire [39:0] _T_562; // @[Frontend.scala 257:34]
  wire  predicted_taken; // @[Frontend.scala 183:29]
  wire [39:0] _T_290; // @[Cat.scala 30:58]
  wire [39:0] _GEN_27; // @[Frontend.scala 183:56]
  wire [39:0] _GEN_42; // @[Frontend.scala 252:61]
  wire [39:0] _GEN_45; // @[Frontend.scala 245:30]
  wire [39:0] _GEN_78; // @[Frontend.scala 252:61]
  wire [39:0] _GEN_81; // @[Frontend.scala 245:30]
  wire [39:0] _GEN_98; // @[Frontend.scala 236:25]
  wire [39:0] predicted_npc; // @[Frontend.scala 296:19]
  wire [39:0] npc; // @[Frontend.scala 120:16]
  wire  _T_252; // @[Frontend.scala 126:53]
  wire  _T_253; // @[Frontend.scala 126:41]
  wire  s0_speculative; // @[Frontend.scala 126:72]
  wire  _T_771; // @[Frontend.scala 221:29]
  wire  _T_772; // @[Frontend.scala 221:53]
  wire  _T_773; // @[Frontend.scala 221:40]
  wire  _T_774; // @[Frontend.scala 221:17]
  wire  _T_642; // @[Frontend.scala 216:26]
  wire  taken_rvcJALR_1; // @[Frontend.scala 216:49]
  wire  _T_775; // @[Frontend.scala 222:27]
  wire  _T_776; // @[Frontend.scala 222:38]
  wire  _T_777; // @[Frontend.scala 222:60]
  wire  _T_778; // @[Frontend.scala 222:47]
  wire  _T_779; // @[Frontend.scala 222:15]
  wire  taken_taken_1; // @[Frontend.scala 221:71]
  wire  taken; // @[Frontend.scala 277:19]
  wire  _GEN_115; // @[Frontend.scala 307:33]
  wire  _GEN_119; // @[Frontend.scala 303:20]
  wire  s2_redirect; // @[Frontend.scala 302:26]
  wire  _GEN_0; // @[Frontend.scala 132:21]
  wire  _T_262; // @[Frontend.scala 153:36]
  wire  _T_265; // @[Frontend.scala 154:39]
  reg  _T_268; // @[Frontend.scala 157:29]
  reg [31:0] _RAND_20;
  wire  _T_269; // @[Frontend.scala 157:40]
  wire  _T_271; // @[Frontend.scala 157:98]
  wire  _T_272; // @[Frontend.scala 157:77]
  wire [39:0] _T_274; // @[Frontend.scala 159:28]
  wire [39:0] _T_276; // @[Frontend.scala 331:33]
  wire [2:0] _T_279; // @[Frontend.scala 162:52]
  wire  _T_281; // @[Frontend.scala 163:76]
  wire  _T_283; // @[Frontend.scala 163:101]
  wire  _T_285; // @[Frontend.scala 167:30]
  wire  fetch_bubble_likely; // @[Frontend.scala 284:33]
  wire  _T_301; // @[Frontend.scala 285:51]
  wire  _T_302; // @[Frontend.scala 285:66]
  wire  _T_841; // @[Frontend.scala 264:52]
  wire  _T_842; // @[Frontend.scala 264:91]
  wire  _T_843; // @[Frontend.scala 264:106]
  wire  _T_844; // @[Frontend.scala 264:34]
  wire  _T_571; // @[Frontend.scala 264:52]
  wire  _T_572; // @[Frontend.scala 264:91]
  wire  _T_573; // @[Frontend.scala 264:106]
  wire  _T_574; // @[Frontend.scala 264:34]
  wire  _GEN_91; // @[Frontend.scala 264:125]
  wire  updateBTB; // @[Frontend.scala 236:25]
  wire  _T_303; // @[Frontend.scala 285:89]
  wire [1:0] _T_304; // @[Frontend.scala 289:63]
  wire [39:0] _GEN_128; // @[Frontend.scala 289:50]
  wire [39:0] _T_305; // @[Frontend.scala 289:50]
  wire [39:0] _GEN_35; // @[Frontend.scala 283:37]
  wire [39:0] _GEN_36; // @[Frontend.scala 283:37]
  wire [1:0] after_idx; // @[Frontend.scala 236:25]
  wire [2:0] _T_306; // @[Frontend.scala 293:66]
  wire [39:0] _GEN_129; // @[Frontend.scala 293:53]
  wire [39:0] _T_308; // @[Frontend.scala 293:53]
  wire  _T_324; // @[Frontend.scala 209:30]
  wire  taken_rviCall; // @[Frontend.scala 209:42]
  wire  _T_521; // @[Frontend.scala 227:22]
  wire  _T_523; // @[Frontend.scala 227:43]
  wire  _T_524; // @[Frontend.scala 227:77]
  wire  _T_526; // @[Frontend.scala 227:86]
  wire  _GEN_38; // @[Frontend.scala 227:95]
  wire  _GEN_39; // @[Frontend.scala 227:95]
  wire  _T_531; // @[Frontend.scala 239:92]
  wire  _T_532; // @[Frontend.scala 239:80]
  wire  _T_533; // @[Frontend.scala 239:127]
  wire  _T_534; // @[Frontend.scala 239:115]
  wire  _T_535; // @[Frontend.scala 239:106]
  wire  _T_536; // @[Frontend.scala 239:68]
  wire  _T_537; // @[Frontend.scala 240:50]
  wire  _T_538; // @[Frontend.scala 241:50]
  wire  _T_539; // @[Frontend.scala 242:50]
  wire  _T_542; // @[Frontend.scala 242:46]
  wire [1:0] _T_543; // @[Frontend.scala 241:46]
  wire [1:0] _T_544; // @[Frontend.scala 240:46]
  wire  _T_547; // @[Frontend.scala 246:34]
  wire  _T_549; // @[Frontend.scala 246:43]
  wire  _T_551; // @[Frontend.scala 246:61]
  wire  _T_553; // @[Frontend.scala 246:77]
  wire  _GEN_40; // @[Frontend.scala 246:96]
  wire  _GEN_43; // @[Frontend.scala 245:30]
  wire  _GEN_46; // @[Frontend.scala 260:59]
  wire  taken_rvc_1; // @[Frontend.scala 199:45]
  wire  _T_591; // @[Frontend.scala 209:30]
  wire  taken_rviCall_1; // @[Frontend.scala 209:42]
  wire  _T_790; // @[Frontend.scala 227:43]
  wire  _T_791; // @[Frontend.scala 227:77]
  wire  _T_793; // @[Frontend.scala 227:86]
  wire  _GEN_75; // @[Frontend.scala 227:95]
  wire  _T_798; // @[Frontend.scala 239:92]
  wire  _T_799; // @[Frontend.scala 239:80]
  wire  _T_800; // @[Frontend.scala 239:127]
  wire  _T_801; // @[Frontend.scala 239:115]
  wire  _T_802; // @[Frontend.scala 239:106]
  wire  _T_803; // @[Frontend.scala 239:68]
  wire  _T_804; // @[Frontend.scala 240:50]
  wire  _T_805; // @[Frontend.scala 241:50]
  wire  _T_806; // @[Frontend.scala 242:50]
  wire  _T_809; // @[Frontend.scala 242:46]
  wire [1:0] _T_810; // @[Frontend.scala 241:46]
  wire [1:0] _T_811; // @[Frontend.scala 240:46]
  wire  _T_814; // @[Frontend.scala 246:34]
  wire  _T_816; // @[Frontend.scala 246:43]
  wire  _T_818; // @[Frontend.scala 246:61]
  wire  _T_820; // @[Frontend.scala 246:77]
  wire  _GEN_76; // @[Frontend.scala 246:96]
  wire  _GEN_82; // @[Frontend.scala 260:59]
  wire  _T_847; // @[Frontend.scala 272:23]
  wire  _T_849; // @[Frontend.scala 272:37]
  wire [15:0] _T_850; // @[Frontend.scala 274:37]
  wire  _T_852; // @[Frontend.scala 299:45]
  wire  _T_853; // @[Frontend.scala 299:28]
  wire  _GEN_116; // @[Frontend.scala 303:20]
  wire  _GEN_117; // @[Frontend.scala 303:20]
  wire [4:0] _GEN_118; // @[Frontend.scala 303:20]
  wire  _T_858; // @[Frontend.scala 311:35]
  wire  _T_860; // @[Frontend.scala 311:11]
  reg [5:0] Frontend_state; // @[Register tracking Frontend state]
  reg [31:0] _RAND_21;
  reg  Frontend_cov [0:63]; // @[Coverage map for Frontend]
  reg [31:0] _RAND_22;
  wire  Frontend_cov_read_data; // @[Coverage map for Frontend]
  wire [5:0] Frontend_cov_read_addr; // @[Coverage map for Frontend]
  wire  Frontend_cov_write_data; // @[Coverage map for Frontend]
  wire [5:0] Frontend_cov_write_addr; // @[Coverage map for Frontend]
  wire  Frontend_cov_write_mask; // @[Coverage map for Frontend]
  wire  Frontend_cov_write_en; // @[Coverage map for Frontend]
  reg [29:0] Frontend_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_23;
  wire  s2_btb_resp_bits_bht_value_shl;
  wire [5:0] s2_btb_resp_bits_bht_value_pad;
  wire [1:0] s2_btb_resp_bits_taken_shl;
  wire [5:0] s2_btb_resp_bits_taken_pad;
  wire [2:0] _T_249_shl;
  wire [5:0] _T_249_pad;
  wire [3:0] s2_partial_insn_valid_shl;
  wire [5:0] s2_partial_insn_valid_pad;
  wire [4:0] s2_btb_resp_valid_shl;
  wire [5:0] s2_btb_resp_valid_pad;
  wire [5:0] s2_valid_shl;
  wire [5:0] s2_valid_pad;
  wire [5:0] Frontend_xor4;
  wire [5:0] Frontend_xor1;
  wire [5:0] Frontend_xor6;
  wire [5:0] Frontend_xor2;
  wire [5:0] Frontend_xor0;
  wire [29:0] icache_sum;
  wire [29:0] fq_sum;
  wire [29:0] tlb_sum;
  wire [29:0] btb_sum;
  wire  stopEn0;
  wire  stopEn1;
  wire  icache_metaAssert_wire;
  wire  fq_metaAssert_wire;
  wire  tlb_metaAssert_wire;
  wire  btb_metaAssert_wire;
  wire  Frontend_or4;
  wire  Frontend_or1;
  wire  Frontend_or6;
  wire  Frontend_or2;
  wire  Frontend_or0;
  ICache icache ( // @[Frontend.scala 61:26]
    .clock(icache_clock),
    .reset(icache_reset),
    .auto_master_out_a_ready(icache_auto_master_out_a_ready),
    .auto_master_out_a_valid(icache_auto_master_out_a_valid),
    .auto_master_out_a_bits_address(icache_auto_master_out_a_bits_address),
    .auto_master_out_d_valid(icache_auto_master_out_d_valid),
    .auto_master_out_d_bits_opcode(icache_auto_master_out_d_bits_opcode),
    .auto_master_out_d_bits_size(icache_auto_master_out_d_bits_size),
    .auto_master_out_d_bits_data(icache_auto_master_out_d_bits_data),
    .auto_master_out_d_bits_corrupt(icache_auto_master_out_d_bits_corrupt),
    .io_req_ready(icache_io_req_ready),
    .io_req_valid(icache_io_req_valid),
    .io_req_bits_addr(icache_io_req_bits_addr),
    .io_s1_paddr(icache_io_s1_paddr),
    .io_s1_kill(icache_io_s1_kill),
    .io_s2_kill(icache_io_s2_kill),
    .io_resp_valid(icache_io_resp_valid),
    .io_resp_bits_data(icache_io_resp_bits_data),
    .io_resp_bits_ae(icache_io_resp_bits_ae),
    .io_invalidate(icache_io_invalidate),
    .io_covSum(icache_io_covSum),
    .metaAssert(icache_metaAssert),
    .metaReset(icache_metaReset)
  );
  ShiftQueue fq ( // @[Frontend.scala 82:57]
    .clock(fq_clock),
    .reset(fq_reset),
    .io_enq_ready(fq_io_enq_ready),
    .io_enq_valid(fq_io_enq_valid),
    .io_enq_bits_btb_taken(fq_io_enq_bits_btb_taken),
    .io_enq_bits_btb_bridx(fq_io_enq_bits_btb_bridx),
    .io_enq_bits_btb_entry(fq_io_enq_bits_btb_entry),
    .io_enq_bits_btb_bht_history(fq_io_enq_bits_btb_bht_history),
    .io_enq_bits_pc(fq_io_enq_bits_pc),
    .io_enq_bits_data(fq_io_enq_bits_data),
    .io_enq_bits_mask(fq_io_enq_bits_mask),
    .io_enq_bits_xcpt_pf_inst(fq_io_enq_bits_xcpt_pf_inst),
    .io_enq_bits_xcpt_ae_inst(fq_io_enq_bits_xcpt_ae_inst),
    .io_enq_bits_replay(fq_io_enq_bits_replay),
    .io_deq_ready(fq_io_deq_ready),
    .io_deq_valid(fq_io_deq_valid),
    .io_deq_bits_btb_taken(fq_io_deq_bits_btb_taken),
    .io_deq_bits_btb_bridx(fq_io_deq_bits_btb_bridx),
    .io_deq_bits_btb_entry(fq_io_deq_bits_btb_entry),
    .io_deq_bits_btb_bht_history(fq_io_deq_bits_btb_bht_history),
    .io_deq_bits_pc(fq_io_deq_bits_pc),
    .io_deq_bits_data(fq_io_deq_bits_data),
    .io_deq_bits_xcpt_pf_inst(fq_io_deq_bits_xcpt_pf_inst),
    .io_deq_bits_xcpt_ae_inst(fq_io_deq_bits_xcpt_ae_inst),
    .io_deq_bits_replay(fq_io_deq_bits_replay),
    .io_mask(fq_io_mask),
    .io_covSum(fq_io_covSum),
    .metaAssert(fq_metaAssert),
    .metaReset(fq_metaReset)
  );
  TLB_1 tlb ( // @[Frontend.scala 95:19]
    .clock(tlb_clock),
    .reset(tlb_reset),
    .io_req_ready(tlb_io_req_ready),
    .io_req_valid(tlb_io_req_valid),
    .io_req_bits_vaddr(tlb_io_req_bits_vaddr),
    .io_resp_miss(tlb_io_resp_miss),
    .io_resp_paddr(tlb_io_resp_paddr),
    .io_resp_pf_inst(tlb_io_resp_pf_inst),
    .io_resp_ae_inst(tlb_io_resp_ae_inst),
    .io_resp_cacheable(tlb_io_resp_cacheable),
    .io_sfence_valid(tlb_io_sfence_valid),
    .io_sfence_bits_rs1(tlb_io_sfence_bits_rs1),
    .io_sfence_bits_rs2(tlb_io_sfence_bits_rs2),
    .io_sfence_bits_addr(tlb_io_sfence_bits_addr),
    .io_ptw_req_ready(tlb_io_ptw_req_ready),
    .io_ptw_req_valid(tlb_io_ptw_req_valid),
    .io_ptw_req_bits_valid(tlb_io_ptw_req_bits_valid),
    .io_ptw_req_bits_bits_addr(tlb_io_ptw_req_bits_bits_addr),
    .io_ptw_resp_valid(tlb_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae(tlb_io_ptw_resp_bits_ae),
    .io_ptw_resp_bits_pte_ppn(tlb_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d(tlb_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(tlb_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(tlb_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(tlb_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(tlb_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(tlb_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(tlb_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(tlb_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(tlb_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous(tlb_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(tlb_io_ptw_ptbr_mode),
    .io_ptw_status_prv(tlb_io_ptw_status_prv),
    .io_ptw_pmp_0_cfg_l(tlb_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a(tlb_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(tlb_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(tlb_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(tlb_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(tlb_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(tlb_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(tlb_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a(tlb_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(tlb_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(tlb_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(tlb_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(tlb_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(tlb_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(tlb_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a(tlb_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(tlb_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(tlb_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(tlb_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(tlb_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(tlb_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(tlb_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a(tlb_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(tlb_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(tlb_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(tlb_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(tlb_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(tlb_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(tlb_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a(tlb_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(tlb_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(tlb_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(tlb_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(tlb_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(tlb_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(tlb_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a(tlb_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(tlb_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(tlb_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(tlb_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(tlb_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(tlb_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(tlb_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a(tlb_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(tlb_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(tlb_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(tlb_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(tlb_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(tlb_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(tlb_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a(tlb_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(tlb_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(tlb_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(tlb_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(tlb_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(tlb_io_ptw_pmp_7_mask),
    .io_ptw_vpoffset_bits_value(tlb_io_ptw_vpoffset_bits_value),
    .io_kill(tlb_io_kill),
    .io_covSum(tlb_io_covSum),
    .metaAssert(tlb_metaAssert),
    .metaReset(tlb_metaReset)
  );
  BTB btb ( // @[Frontend.scala 170:21]
    .clock(btb_clock),
    .reset(btb_reset),
    .io_req_bits_addr(btb_io_req_bits_addr),
    .io_resp_valid(btb_io_resp_valid),
    .io_resp_bits_taken(btb_io_resp_bits_taken),
    .io_resp_bits_bridx(btb_io_resp_bits_bridx),
    .io_resp_bits_target(btb_io_resp_bits_target),
    .io_resp_bits_entry(btb_io_resp_bits_entry),
    .io_resp_bits_bht_history(btb_io_resp_bits_bht_history),
    .io_resp_bits_bht_value(btb_io_resp_bits_bht_value),
    .io_btb_update_valid(btb_io_btb_update_valid),
    .io_btb_update_bits_prediction_entry(btb_io_btb_update_bits_prediction_entry),
    .io_btb_update_bits_pc(btb_io_btb_update_bits_pc),
    .io_btb_update_bits_isValid(btb_io_btb_update_bits_isValid),
    .io_btb_update_bits_br_pc(btb_io_btb_update_bits_br_pc),
    .io_btb_update_bits_cfiType(btb_io_btb_update_bits_cfiType),
    .io_bht_update_valid(btb_io_bht_update_valid),
    .io_bht_update_bits_prediction_history(btb_io_bht_update_bits_prediction_history),
    .io_bht_update_bits_pc(btb_io_bht_update_bits_pc),
    .io_bht_update_bits_branch(btb_io_bht_update_bits_branch),
    .io_bht_update_bits_taken(btb_io_bht_update_bits_taken),
    .io_bht_update_bits_mispredict(btb_io_bht_update_bits_mispredict),
    .io_bht_advance_valid(btb_io_bht_advance_valid),
    .io_bht_advance_bits_bht_value(btb_io_bht_advance_bits_bht_value),
    .io_ras_update_valid(btb_io_ras_update_valid),
    .io_ras_update_bits_cfiType(btb_io_ras_update_bits_cfiType),
    .io_ras_update_bits_returnAddr(btb_io_ras_update_bits_returnAddr),
    .io_ras_head_valid(btb_io_ras_head_valid),
    .io_ras_head_bits(btb_io_ras_head_bits),
    .io_flush(btb_io_flush),
    .io_covSum(btb_io_covSum),
    .metaAssert(btb_metaAssert),
    .metaReset(btb_metaReset)
  );
  assign _T_212 = io_cpu_req_valid | io_cpu_sfence_valid; // @[Frontend.scala 86:29]
  assign _T_213 = _T_212 | io_cpu_flush_icache; // @[Frontend.scala 86:52]
  assign _T_214 = _T_213 | io_cpu_bht_update_valid; // @[Frontend.scala 86:75]
  assign _T_215 = _T_214 | io_cpu_btb_update_valid; // @[Frontend.scala 86:102]
  assign _T_217 = ~_T_215 | io_cpu_might_request; // @[Frontend.scala 86:130]
  assign _T_219 = _T_217 | reset; // @[Frontend.scala 86:9]
  assign s0_valid = io_cpu_req_valid | ~fq_io_mask[2]; // @[Frontend.scala 97:35]
  assign _T_229 = ~io_reset_vector | 32'h1; // @[Frontend.scala 331:33]
  assign s2_btb_taken = s2_btb_resp_valid & s2_btb_resp_bits_taken; // @[Frontend.scala 105:40]
  assign s2_xcpt = s2_tlb_resp_ae_inst | s2_tlb_resp_pf_inst; // @[Frontend.scala 107:37]
  assign _T_238 = ~s1_pc | 40'h3; // @[Frontend.scala 113:29]
  assign s1_base_pc = ~_T_238; // @[Frontend.scala 113:20]
  assign ntpc = s1_base_pc + 40'h4; // @[Frontend.scala 114:25]
  assign _T_243 = fq_io_enq_ready & fq_io_enq_valid; // @[Decoupled.scala 37:37]
  assign _T_245 = s2_valid & ~_T_243; // @[Frontend.scala 119:26]
  assign s2_replay = _T_245 | _T_249; // @[Frontend.scala 119:48]
  assign _T_247 = s2_replay & ~s0_valid; // @[Frontend.scala 119:69]
  assign _T_310 = s2_partial_insn[1:0] != 2'h3; // @[Frontend.scala 199:45]
  assign taken_prevRVI = s2_partial_insn_valid & ~_T_310; // @[Frontend.scala 200:31]
  assign taken_bits = fq_io_enq_bits_data[15:0]; // @[Frontend.scala 202:37]
  assign taken_rviBits = {taken_bits,s2_partial_insn}; // @[Cat.scala 30:58]
  assign taken_rviJump = taken_rviBits[6:0] == 7'h6f; // @[Frontend.scala 206:34]
  assign taken_rviJALR = taken_rviBits[6:0] == 7'h67; // @[Frontend.scala 207:34]
  assign _T_504 = taken_rviJump | taken_rviJALR; // @[Frontend.scala 221:29]
  assign taken_rviBranch = taken_rviBits[6:0] == 7'h63; // @[Frontend.scala 205:36]
  assign _T_505 = taken_rviBranch & s2_btb_resp_bits_bht_value; // @[Frontend.scala 221:53]
  assign _T_506 = _T_504 | _T_505; // @[Frontend.scala 221:40]
  assign _T_507 = taken_prevRVI & _T_506; // @[Frontend.scala 221:17]
  assign taken_valid = fq_io_enq_bits_mask[0] & ~taken_prevRVI; // @[Frontend.scala 201:44]
  assign _T_332 = taken_bits & 16'he003; // @[Frontend.scala 212:26]
  assign taken_rvcJump = 16'ha001 == _T_332; // @[Frontend.scala 212:26]
  assign _T_374 = taken_bits & 16'hf003; // @[Frontend.scala 216:26]
  assign _T_375 = 16'h9002 == _T_374; // @[Frontend.scala 216:26]
  assign _T_377 = taken_bits[6:2] == 5'h0; // @[Frontend.scala 216:62]
  assign taken_rvcJALR = _T_375 & _T_377; // @[Frontend.scala 216:49]
  assign _T_508 = taken_rvcJump | taken_rvcJALR; // @[Frontend.scala 222:27]
  assign _T_368 = 16'h8002 == _T_374; // @[Frontend.scala 214:24]
  assign taken_rvcJR = _T_368 & _T_377; // @[Frontend.scala 214:46]
  assign _T_509 = _T_508 | taken_rvcJR; // @[Frontend.scala 222:38]
  assign _T_327 = 16'hc001 == _T_332; // @[Frontend.scala 210:28]
  assign _T_329 = 16'he001 == _T_332; // @[Frontend.scala 210:60]
  assign taken_rvcBranch = _T_327 | _T_329; // @[Frontend.scala 210:52]
  assign _T_510 = taken_rvcBranch & s2_btb_resp_bits_bht_value; // @[Frontend.scala 222:60]
  assign _T_511 = _T_509 | _T_510; // @[Frontend.scala 222:47]
  assign _T_512 = taken_valid & _T_511; // @[Frontend.scala 222:15]
  assign taken_taken = _T_507 | _T_512; // @[Frontend.scala 221:71]
  assign taken_idx = ~taken_taken; // @[Frontend.scala 236:13]
  assign _T_577 = taken_bits[1:0] != 2'h3; // @[Frontend.scala 199:45]
  assign taken_prevRVI_1 = taken_valid & ~_T_577; // @[Frontend.scala 200:31]
  assign taken_bits_1 = fq_io_enq_bits_data[31:16]; // @[Frontend.scala 202:37]
  assign taken_rviBits_1 = {taken_bits_1,taken_bits}; // @[Cat.scala 30:58]
  assign taken_rviJALR_1 = taken_rviBits_1[6:0] == 7'h67; // @[Frontend.scala 207:34]
  assign _T_587 = taken_rviJALR_1 & ~taken_rviBits_1[7]; // @[Frontend.scala 208:31]
  assign _T_589 = taken_rviBits_1[19:15] & 5'h1b; // @[Frontend.scala 208:66]
  assign _T_590 = 5'h1 == _T_589; // @[Frontend.scala 208:66]
  assign taken_rviReturn_1 = _T_587 & _T_590; // @[Frontend.scala 208:46]
  assign _T_780 = taken_prevRVI_1 & taken_rviReturn_1; // @[Frontend.scala 223:61]
  assign taken_valid_1 = fq_io_enq_bits_mask[1] & ~taken_prevRVI_1; // @[Frontend.scala 201:44]
  assign _T_634 = taken_bits_1 & 16'hf003; // @[Frontend.scala 214:24]
  assign _T_635 = 16'h8002 == _T_634; // @[Frontend.scala 214:24]
  assign _T_637 = taken_bits_1[6:2] == 5'h0; // @[Frontend.scala 214:59]
  assign taken_rvcJR_1 = _T_635 & _T_637; // @[Frontend.scala 214:46]
  assign _T_639 = taken_bits_1[11:7] & 5'h1b; // @[Frontend.scala 215:49]
  assign _T_640 = 5'h1 == _T_639; // @[Frontend.scala 215:49]
  assign taken_rvcReturn_1 = taken_rvcJR_1 & _T_640; // @[Frontend.scala 215:29]
  assign _T_781 = taken_valid_1 & taken_rvcReturn_1; // @[Frontend.scala 223:83]
  assign _T_782 = _T_780 | _T_781; // @[Frontend.scala 223:74]
  assign taken_predictReturn_1 = btb_io_ras_head_valid & _T_782; // @[Frontend.scala 223:49]
  assign _T_821 = s2_valid & taken_predictReturn_1; // @[Frontend.scala 249:26]
  assign _T_320 = taken_rviJALR & ~taken_rviBits[7]; // @[Frontend.scala 208:31]
  assign _T_322 = taken_rviBits[19:15] & 5'h1b; // @[Frontend.scala 208:66]
  assign _T_323 = 5'h1 == _T_322; // @[Frontend.scala 208:66]
  assign taken_rviReturn = _T_320 & _T_323; // @[Frontend.scala 208:46]
  assign _T_513 = taken_prevRVI & taken_rviReturn; // @[Frontend.scala 223:61]
  assign _T_372 = taken_bits[11:7] & 5'h1b; // @[Frontend.scala 215:49]
  assign _T_373 = 5'h1 == _T_372; // @[Frontend.scala 215:49]
  assign taken_rvcReturn = taken_rvcJR & _T_373; // @[Frontend.scala 215:29]
  assign _T_514 = taken_valid & taken_rvcReturn; // @[Frontend.scala 223:83]
  assign _T_515 = _T_513 | _T_514; // @[Frontend.scala 223:74]
  assign taken_predictReturn = btb_io_ras_head_valid & _T_515; // @[Frontend.scala 223:49]
  assign _T_554 = s2_valid & taken_predictReturn; // @[Frontend.scala 249:26]
  assign _GEN_44 = ~s2_btb_taken & _T_554; // @[Frontend.scala 245:30]
  assign _GEN_77 = _T_821 | _GEN_44; // @[Frontend.scala 249:44]
  assign _GEN_80 = s2_btb_taken ? _GEN_44 : _GEN_77; // @[Frontend.scala 245:30]
  assign useRAS = taken_idx ? _GEN_80 : _GEN_44; // @[Frontend.scala 236:25]
  assign taken_rviBranch_1 = taken_rviBits_1[6:0] == 7'h63; // @[Frontend.scala 205:36]
  assign _T_785 = taken_prevRVI_1 & taken_rviBranch_1; // @[Frontend.scala 225:53]
  assign _T_593 = taken_bits_1 & 16'he003; // @[Frontend.scala 210:28]
  assign _T_594 = 16'hc001 == _T_593; // @[Frontend.scala 210:28]
  assign _T_596 = 16'he001 == _T_593; // @[Frontend.scala 210:60]
  assign taken_rvcBranch_1 = _T_594 | _T_596; // @[Frontend.scala 210:52]
  assign _T_786 = taken_valid_1 & taken_rvcBranch_1; // @[Frontend.scala 225:75]
  assign _T_787 = _T_785 | _T_786; // @[Frontend.scala 225:66]
  assign taken_predictBranch_1 = s2_btb_resp_bits_bht_value & _T_787; // @[Frontend.scala 225:41]
  assign taken_rviJump_1 = taken_rviBits_1[6:0] == 7'h6f; // @[Frontend.scala 206:34]
  assign _T_783 = taken_prevRVI_1 & taken_rviJump_1; // @[Frontend.scala 224:33]
  assign taken_rvcJump_1 = 16'ha001 == _T_593; // @[Frontend.scala 212:26]
  assign _T_784 = taken_valid_1 & taken_rvcJump_1; // @[Frontend.scala 224:53]
  assign taken_predictJump_1 = _T_783 | _T_784; // @[Frontend.scala 224:44]
  assign _T_822 = taken_predictBranch_1 | taken_predictJump_1; // @[Frontend.scala 252:44]
  assign _T_823 = s2_valid & _T_822; // @[Frontend.scala 252:26]
  assign _T_292 = ~s2_pc | 40'h3; // @[Frontend.scala 192:31]
  assign s2_base_pc = ~_T_292; // @[Frontend.scala 192:22]
  assign taken_pc_1 = s2_base_pc | 40'h2; // @[Frontend.scala 253:33]
  assign _T_826 = taken_pc_1 - 40'h2; // @[Frontend.scala 256:36]
  assign _T_828 = taken_prevRVI_1 ? _T_826 : taken_pc_1; // @[Frontend.scala 256:57]
  assign _T_648 = taken_rviBits_1[31]; // @[RocketCore.scala 954:53]
  assign _T_703 = taken_rviBits_1[31]; // @[Cat.scala 30:58]
  assign _T_702 = {11{_T_648}}; // @[Cat.scala 30:58]
  assign _T_700 = taken_rviBits_1[19:12]; // @[Cat.scala 30:58]
  assign _T_699 = taken_rviBits_1[20]; // @[Cat.scala 30:58]
  assign _T_707 = {_T_703,_T_702,_T_700,_T_699,taken_rviBits_1[30:25],taken_rviBits_1[24:21],1'h0}; // @[RocketCore.scala 968:53]
  assign _T_762 = {8{_T_648}}; // @[Cat.scala 30:58]
  assign _T_761 = taken_rviBits_1[7]; // @[Cat.scala 30:58]
  assign _T_769 = {_T_703,_T_702,_T_762,_T_761,taken_rviBits_1[30:25],taken_rviBits_1[11:8],1'h0}; // @[RocketCore.scala 968:53]
  assign taken_rviImm_1 = taken_rviBits_1[3] ? $signed(_T_707) : $signed(_T_769); // @[Frontend.scala 218:23]
  assign _T_604 = taken_bits_1[12] ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12]
  assign _T_614 = {_T_604,taken_bits_1[6:5],taken_bits_1[2],taken_bits_1[11:10],taken_bits_1[4:3],1'h0}; // @[Frontend.scala 213:66]
  assign _T_617 = taken_bits_1[12] ? 10'h3ff : 10'h0; // @[Bitwise.scala 72:12]
  assign _T_633 = {_T_617,taken_bits_1[8],taken_bits_1[10:9],taken_bits_1[6],taken_bits_1[7],taken_bits_1[2],taken_bits_1[11],taken_bits_1[5:3],1'h0}; // @[Frontend.scala 213:106]
  assign taken_rvcImm_1 = taken_bits_1[14] ? $signed({{8{_T_614[12]}},_T_614}) : $signed(_T_633); // @[Frontend.scala 213:23]
  assign _T_829 = taken_prevRVI_1 ? $signed(taken_rviImm_1) : $signed({{11{taken_rvcImm_1[20]}},taken_rvcImm_1}); // @[Frontend.scala 256:69]
  assign _GEN_126 = {{8{_T_829[31]}},_T_829}; // @[Frontend.scala 256:64]
  assign _T_832 = $signed(_T_828) + $signed(_GEN_126); // @[Frontend.scala 257:34]
  assign _T_518 = taken_prevRVI & taken_rviBranch; // @[Frontend.scala 225:53]
  assign _T_519 = taken_valid & taken_rvcBranch; // @[Frontend.scala 225:75]
  assign _T_520 = _T_518 | _T_519; // @[Frontend.scala 225:66]
  assign taken_predictBranch = s2_btb_resp_bits_bht_value & _T_520; // @[Frontend.scala 225:41]
  assign _T_516 = taken_prevRVI & taken_rviJump; // @[Frontend.scala 224:33]
  assign _T_517 = taken_valid & taken_rvcJump; // @[Frontend.scala 224:53]
  assign taken_predictJump = _T_516 | _T_517; // @[Frontend.scala 224:44]
  assign _T_555 = taken_predictBranch | taken_predictJump; // @[Frontend.scala 252:44]
  assign _T_556 = s2_valid & _T_555; // @[Frontend.scala 252:26]
  assign _T_557 = ~_T_292; // @[Frontend.scala 255:32]
  assign _T_381 = taken_rviBits[31]; // @[RocketCore.scala 954:53]
  assign _T_436 = taken_rviBits[31]; // @[Cat.scala 30:58]
  assign _T_435 = {11{_T_381}}; // @[Cat.scala 30:58]
  assign _T_433 = taken_rviBits[19:12]; // @[Cat.scala 30:58]
  assign _T_432 = taken_rviBits[20]; // @[Cat.scala 30:58]
  assign _T_440 = {_T_436,_T_435,_T_433,_T_432,taken_rviBits[30:25],taken_rviBits[24:21],1'h0}; // @[RocketCore.scala 968:53]
  assign _T_495 = {8{_T_381}}; // @[Cat.scala 30:58]
  assign _T_494 = taken_rviBits[7]; // @[Cat.scala 30:58]
  assign _T_502 = {_T_436,_T_435,_T_495,_T_494,taken_rviBits[30:25],taken_rviBits[11:8],1'h0}; // @[RocketCore.scala 968:53]
  assign taken_rviImm = taken_rviBits[3] ? $signed(_T_440) : $signed(_T_502); // @[Frontend.scala 218:23]
  assign _T_558 = $signed(taken_rviImm) - 32'sh2; // @[Frontend.scala 255:61]
  assign _T_337 = taken_bits[12] ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12]
  assign _T_347 = {_T_337,taken_bits[6:5],taken_bits[2],taken_bits[11:10],taken_bits[4:3],1'h0}; // @[Frontend.scala 213:66]
  assign _T_350 = taken_bits[12] ? 10'h3ff : 10'h0; // @[Bitwise.scala 72:12]
  assign _T_366 = {_T_350,taken_bits[8],taken_bits[10:9],taken_bits[6],taken_bits[7],taken_bits[2],taken_bits[11],taken_bits[5:3],1'h0}; // @[Frontend.scala 213:106]
  assign taken_rvcImm = taken_bits[14] ? $signed({{8{_T_347[12]}},_T_347}) : $signed(_T_366); // @[Frontend.scala 213:23]
  assign _T_559 = taken_prevRVI ? $signed(_T_558) : $signed({{12{taken_rvcImm[20]}},taken_rvcImm}); // @[Frontend.scala 255:44]
  assign _GEN_127 = {{7{_T_559[32]}},_T_559}; // @[Frontend.scala 255:39]
  assign _T_562 = $signed(_T_557) + $signed(_GEN_127); // @[Frontend.scala 257:34]
  assign predicted_taken = btb_io_resp_valid & btb_io_resp_bits_taken; // @[Frontend.scala 183:29]
  assign _T_290 = {btb_io_resp_bits_target[38],btb_io_resp_bits_target}; // @[Cat.scala 30:58]
  assign _GEN_27 = predicted_taken ? _T_290 : ntpc; // @[Frontend.scala 183:56]
  assign _GEN_42 = _T_556 ? _T_562 : _GEN_27; // @[Frontend.scala 252:61]
  assign _GEN_45 = s2_btb_taken ? _GEN_27 : _GEN_42; // @[Frontend.scala 245:30]
  assign _GEN_78 = _T_823 ? _T_832 : _GEN_45; // @[Frontend.scala 252:61]
  assign _GEN_81 = s2_btb_taken ? _GEN_45 : _GEN_78; // @[Frontend.scala 245:30]
  assign _GEN_98 = taken_idx ? _GEN_81 : _GEN_45; // @[Frontend.scala 236:25]
  assign predicted_npc = useRAS ? {{1'd0}, btb_io_ras_head_bits} : _GEN_98; // @[Frontend.scala 296:19]
  assign npc = s2_replay ? s2_pc : predicted_npc; // @[Frontend.scala 120:16]
  assign _T_252 = s2_valid & ~s2_speculative; // @[Frontend.scala 126:53]
  assign _T_253 = s1_speculative | _T_252; // @[Frontend.scala 126:41]
  assign s0_speculative = _T_253 | predicted_taken; // @[Frontend.scala 126:72]
  assign _T_771 = taken_rviJump_1 | taken_rviJALR_1; // @[Frontend.scala 221:29]
  assign _T_772 = taken_rviBranch_1 & s2_btb_resp_bits_bht_value; // @[Frontend.scala 221:53]
  assign _T_773 = _T_771 | _T_772; // @[Frontend.scala 221:40]
  assign _T_774 = taken_prevRVI_1 & _T_773; // @[Frontend.scala 221:17]
  assign _T_642 = 16'h9002 == _T_634; // @[Frontend.scala 216:26]
  assign taken_rvcJALR_1 = _T_642 & _T_637; // @[Frontend.scala 216:49]
  assign _T_775 = taken_rvcJump_1 | taken_rvcJALR_1; // @[Frontend.scala 222:27]
  assign _T_776 = _T_775 | taken_rvcJR_1; // @[Frontend.scala 222:38]
  assign _T_777 = taken_rvcBranch_1 & s2_btb_resp_bits_bht_value; // @[Frontend.scala 222:60]
  assign _T_778 = _T_776 | _T_777; // @[Frontend.scala 222:47]
  assign _T_779 = taken_valid_1 & _T_778; // @[Frontend.scala 222:15]
  assign taken_taken_1 = _T_774 | _T_779; // @[Frontend.scala 221:71]
  assign taken = taken_taken | taken_taken_1; // @[Frontend.scala 277:19]
  assign _GEN_115 = _T_243 | io_cpu_req_valid; // @[Frontend.scala 307:33]
  assign _GEN_119 = taken ? _GEN_115 : io_cpu_req_valid; // @[Frontend.scala 303:20]
  assign s2_redirect = s2_btb_taken ? io_cpu_req_valid : _GEN_119; // @[Frontend.scala 302:26]
  assign _GEN_0 = ~s2_replay & ~s2_redirect; // @[Frontend.scala 132:21]
  assign _T_262 = s2_redirect | tlb_io_resp_miss; // @[Frontend.scala 153:36]
  assign _T_265 = s2_speculative & ~s2_tlb_resp_cacheable; // @[Frontend.scala 154:39]
  assign _T_269 = _T_268 & s2_valid; // @[Frontend.scala 157:40]
  assign _T_271 = ~s2_tlb_resp_miss & icache_io_s2_kill; // @[Frontend.scala 157:98]
  assign _T_272 = icache_io_resp_valid | _T_271; // @[Frontend.scala 157:77]
  assign _T_274 = io_cpu_req_valid ? io_cpu_req_bits_pc : npc; // @[Frontend.scala 159:28]
  assign _T_276 = ~_T_274 | 40'h1; // @[Frontend.scala 331:33]
  assign _T_279 = 3'h3 << s2_pc[1]; // @[Frontend.scala 162:52]
  assign _T_281 = icache_io_s2_kill & ~icache_io_resp_valid; // @[Frontend.scala 163:76]
  assign _T_283 = _T_281 & ~s2_xcpt; // @[Frontend.scala 163:101]
  assign _T_285 = icache_io_resp_valid & icache_io_resp_bits_ae; // @[Frontend.scala 167:30]
  assign fetch_bubble_likely = ~fq_io_mask[1]; // @[Frontend.scala 284:33]
  assign _T_301 = _T_243 & ~wrong_path; // @[Frontend.scala 285:51]
  assign _T_302 = _T_301 & fetch_bubble_likely; // @[Frontend.scala 285:66]
  assign _T_841 = taken_predictBranch_1 & s2_btb_resp_bits_bht_value; // @[Frontend.scala 264:52]
  assign _T_842 = _T_841 | taken_predictJump_1; // @[Frontend.scala 264:91]
  assign _T_843 = _T_842 | taken_predictReturn_1; // @[Frontend.scala 264:106]
  assign _T_844 = ~s2_btb_resp_valid & _T_843; // @[Frontend.scala 264:34]
  assign _T_571 = taken_predictBranch & s2_btb_resp_bits_bht_value; // @[Frontend.scala 264:52]
  assign _T_572 = _T_571 | taken_predictJump; // @[Frontend.scala 264:91]
  assign _T_573 = _T_572 | taken_predictReturn; // @[Frontend.scala 264:106]
  assign _T_574 = ~s2_btb_resp_valid & _T_573; // @[Frontend.scala 264:34]
  assign _GEN_91 = _T_844 | _T_574; // @[Frontend.scala 264:125]
  assign updateBTB = taken_idx ? _GEN_91 : _T_574; // @[Frontend.scala 236:25]
  assign _T_303 = _T_302 & updateBTB; // @[Frontend.scala 285:89]
  assign _T_304 = {taken_idx, 1'h0}; // @[Frontend.scala 289:63]
  assign _GEN_128 = {{38'd0}, _T_304}; // @[Frontend.scala 289:50]
  assign _T_305 = s2_base_pc | _GEN_128; // @[Frontend.scala 289:50]
  assign _GEN_35 = io_cpu_btb_update_valid ? {{1'd0}, io_cpu_btb_update_bits_br_pc} : _T_305; // @[Frontend.scala 283:37]
  assign _GEN_36 = io_cpu_btb_update_valid ? {{1'd0}, io_cpu_btb_update_bits_pc} : s2_base_pc; // @[Frontend.scala 283:37]
  assign after_idx = taken_idx ? 2'h2 : 2'h1; // @[Frontend.scala 236:25]
  assign _T_306 = {after_idx, 1'h0}; // @[Frontend.scala 293:66]
  assign _GEN_129 = {{37'd0}, _T_306}; // @[Frontend.scala 293:53]
  assign _T_308 = s2_base_pc + _GEN_129; // @[Frontend.scala 293:53]
  assign _T_324 = taken_rviJALR | taken_rviJump; // @[Frontend.scala 209:30]
  assign taken_rviCall = _T_324 & taken_rviBits[7]; // @[Frontend.scala 209:42]
  assign _T_521 = s2_valid & s2_btb_resp_valid; // @[Frontend.scala 227:22]
  assign _T_523 = _T_521 & ~s2_btb_resp_bits_bridx; // @[Frontend.scala 227:43]
  assign _T_524 = _T_523 & taken_valid; // @[Frontend.scala 227:77]
  assign _T_526 = _T_524 & ~_T_577; // @[Frontend.scala 227:86]
  assign _GEN_38 = _T_526 | _T_283; // @[Frontend.scala 227:95]
  assign _GEN_39 = _T_526 | wrong_path; // @[Frontend.scala 227:95]
  assign _T_531 = taken_rviCall | taken_rviReturn; // @[Frontend.scala 239:92]
  assign _T_532 = taken_prevRVI & _T_531; // @[Frontend.scala 239:80]
  assign _T_533 = taken_rvcJALR | taken_rvcReturn; // @[Frontend.scala 239:127]
  assign _T_534 = taken_valid & _T_533; // @[Frontend.scala 239:115]
  assign _T_535 = _T_532 | _T_534; // @[Frontend.scala 239:106]
  assign _T_536 = _T_301 & _T_535; // @[Frontend.scala 239:68]
  assign _T_537 = taken_prevRVI ? taken_rviReturn : taken_rvcReturn; // @[Frontend.scala 240:50]
  assign _T_538 = taken_prevRVI ? taken_rviCall : taken_rvcJALR; // @[Frontend.scala 241:50]
  assign _T_539 = taken_prevRVI ? taken_rviBranch : taken_rvcBranch; // @[Frontend.scala 242:50]
  assign _T_542 = _T_539 ? 1'h0 : 1'h1; // @[Frontend.scala 242:46]
  assign _T_543 = _T_538 ? 2'h2 : {{1'd0}, _T_542}; // @[Frontend.scala 241:46]
  assign _T_544 = _T_537 ? 2'h3 : _T_543; // @[Frontend.scala 240:46]
  assign _T_547 = _T_243 & taken_taken; // @[Frontend.scala 246:34]
  assign _T_549 = _T_547 & ~taken_predictBranch; // @[Frontend.scala 246:43]
  assign _T_551 = _T_549 & ~taken_predictJump; // @[Frontend.scala 246:61]
  assign _T_553 = _T_551 & ~taken_predictReturn; // @[Frontend.scala 246:77]
  assign _GEN_40 = _T_553 | _GEN_39; // @[Frontend.scala 246:96]
  assign _GEN_43 = s2_btb_taken ? _GEN_39 : _GEN_40; // @[Frontend.scala 245:30]
  assign _GEN_46 = _T_520 & _T_301; // @[Frontend.scala 260:59]
  assign taken_rvc_1 = taken_bits_1[1:0] != 2'h3; // @[Frontend.scala 199:45]
  assign _T_591 = taken_rviJALR_1 | taken_rviJump_1; // @[Frontend.scala 209:30]
  assign taken_rviCall_1 = _T_591 & taken_rviBits_1[7]; // @[Frontend.scala 209:42]
  assign _T_790 = _T_521 & s2_btb_resp_bits_bridx; // @[Frontend.scala 227:43]
  assign _T_791 = _T_790 & taken_valid_1; // @[Frontend.scala 227:77]
  assign _T_793 = _T_791 & ~taken_rvc_1; // @[Frontend.scala 227:86]
  assign _GEN_75 = _T_793 | _GEN_43; // @[Frontend.scala 227:95]
  assign _T_798 = taken_rviCall_1 | taken_rviReturn_1; // @[Frontend.scala 239:92]
  assign _T_799 = taken_prevRVI_1 & _T_798; // @[Frontend.scala 239:80]
  assign _T_800 = taken_rvcJALR_1 | taken_rvcReturn_1; // @[Frontend.scala 239:127]
  assign _T_801 = taken_valid_1 & _T_800; // @[Frontend.scala 239:115]
  assign _T_802 = _T_799 | _T_801; // @[Frontend.scala 239:106]
  assign _T_803 = _T_301 & _T_802; // @[Frontend.scala 239:68]
  assign _T_804 = taken_prevRVI_1 ? taken_rviReturn_1 : taken_rvcReturn_1; // @[Frontend.scala 240:50]
  assign _T_805 = taken_prevRVI_1 ? taken_rviCall_1 : taken_rvcJALR_1; // @[Frontend.scala 241:50]
  assign _T_806 = taken_prevRVI_1 ? taken_rviBranch_1 : taken_rvcBranch_1; // @[Frontend.scala 242:50]
  assign _T_809 = _T_806 ? 1'h0 : 1'h1; // @[Frontend.scala 242:46]
  assign _T_810 = _T_805 ? 2'h2 : {{1'd0}, _T_809}; // @[Frontend.scala 241:46]
  assign _T_811 = _T_804 ? 2'h3 : _T_810; // @[Frontend.scala 240:46]
  assign _T_814 = _T_243 & taken_taken_1; // @[Frontend.scala 246:34]
  assign _T_816 = _T_814 & ~taken_predictBranch_1; // @[Frontend.scala 246:43]
  assign _T_818 = _T_816 & ~taken_predictJump_1; // @[Frontend.scala 246:61]
  assign _T_820 = _T_818 & ~taken_predictReturn_1; // @[Frontend.scala 246:77]
  assign _GEN_76 = _T_820 | _GEN_75; // @[Frontend.scala 246:96]
  assign _GEN_82 = _T_787 ? _T_301 : _GEN_46; // @[Frontend.scala 260:59]
  assign _T_847 = taken_valid_1 & taken_idx; // @[Frontend.scala 272:23]
  assign _T_849 = _T_847 & ~taken_rvc_1; // @[Frontend.scala 272:37]
  assign _T_850 = taken_bits_1 | 16'h3; // @[Frontend.scala 274:37]
  assign _T_852 = s2_btb_taken | taken; // @[Frontend.scala 299:45]
  assign _T_853 = _T_243 & _T_852; // @[Frontend.scala 299:28]
  assign _GEN_116 = taken ? taken_idx : s2_btb_resp_bits_bridx; // @[Frontend.scala 303:20]
  assign _GEN_117 = taken | s2_btb_taken; // @[Frontend.scala 303:20]
  assign _GEN_118 = taken ? 5'h1c : s2_btb_resp_bits_entry; // @[Frontend.scala 303:20]
  assign _T_858 = ~s2_partial_insn_valid | fq_io_enq_bits_mask[0]; // @[Frontend.scala 311:35]
  assign _T_860 = _T_858 | reset; // @[Frontend.scala 311:11]
  assign auto_icache_master_out_a_valid = icache_auto_master_out_a_valid; // @[LazyModule.scala 173:49]
  assign auto_icache_master_out_a_bits_address = icache_auto_master_out_a_bits_address; // @[LazyModule.scala 173:49]
  assign io_cpu_resp_valid = fq_io_deq_valid; // @[Frontend.scala 316:15]
  assign io_cpu_resp_bits_btb_taken = fq_io_deq_bits_btb_taken; // @[Frontend.scala 316:15]
  assign io_cpu_resp_bits_btb_bridx = fq_io_deq_bits_btb_bridx; // @[Frontend.scala 316:15]
  assign io_cpu_resp_bits_btb_entry = fq_io_deq_bits_btb_entry; // @[Frontend.scala 316:15]
  assign io_cpu_resp_bits_btb_bht_history = fq_io_deq_bits_btb_bht_history; // @[Frontend.scala 316:15]
  assign io_cpu_resp_bits_pc = fq_io_deq_bits_pc; // @[Frontend.scala 316:15]
  assign io_cpu_resp_bits_data = fq_io_deq_bits_data; // @[Frontend.scala 316:15]
  assign io_cpu_resp_bits_xcpt_pf_inst = fq_io_deq_bits_xcpt_pf_inst; // @[Frontend.scala 316:15]
  assign io_cpu_resp_bits_xcpt_ae_inst = fq_io_deq_bits_xcpt_ae_inst; // @[Frontend.scala 316:15]
  assign io_cpu_resp_bits_replay = fq_io_deq_bits_replay; // @[Frontend.scala 316:15]
  assign io_cpu_npc = ~_T_276; // @[Frontend.scala 159:14]
  assign io_ptw_req_valid = tlb_io_ptw_req_valid; // @[Frontend.scala 139:10]
  assign io_ptw_req_bits_valid = tlb_io_ptw_req_bits_valid; // @[Frontend.scala 139:10]
  assign io_ptw_req_bits_bits_addr = tlb_io_ptw_req_bits_bits_addr; // @[Frontend.scala 139:10]
  assign icache_clock = gated_clock; // @[Frontend.scala 91:16]
  assign icache_reset = reset;
  assign icache_auto_master_out_a_ready = auto_icache_master_out_a_ready; // @[LazyModule.scala 173:49]
  assign icache_auto_master_out_d_valid = auto_icache_master_out_d_valid; // @[LazyModule.scala 173:49]
  assign icache_auto_master_out_d_bits_opcode = auto_icache_master_out_d_bits_opcode; // @[LazyModule.scala 173:49]
  assign icache_auto_master_out_d_bits_size = auto_icache_master_out_d_bits_size; // @[LazyModule.scala 173:49]
  assign icache_auto_master_out_d_bits_data = auto_icache_master_out_d_bits_data; // @[LazyModule.scala 173:49]
  assign icache_auto_master_out_d_bits_corrupt = auto_icache_master_out_d_bits_corrupt; // @[LazyModule.scala 173:49]
  assign icache_io_req_valid = io_cpu_req_valid | ~fq_io_mask[2]; // @[Frontend.scala 148:23]
  assign icache_io_req_bits_addr = io_cpu_npc[38:0]; // @[Frontend.scala 149:27]
  assign icache_io_s1_paddr = tlb_io_resp_paddr; // @[Frontend.scala 151:22]
  assign icache_io_s1_kill = _T_262 | s2_replay; // @[Frontend.scala 153:21]
  assign icache_io_s2_kill = _T_265 | s2_xcpt; // @[Frontend.scala 154:21]
  assign icache_io_invalidate = io_cpu_flush_icache; // @[Frontend.scala 150:24]
  assign fq_clock = gated_clock;
  assign fq_reset = reset | io_cpu_req_valid;
  assign fq_io_enq_valid = _T_269 & _T_272; // @[Frontend.scala 157:19]
  assign fq_io_enq_bits_btb_taken = s2_btb_taken ? s2_btb_taken : _GEN_117; // @[Frontend.scala 164:22 Frontend.scala 165:28 Frontend.scala 305:34]
  assign fq_io_enq_bits_btb_bridx = s2_btb_taken ? s2_btb_resp_bits_bridx : _GEN_116; // @[Frontend.scala 164:22 Frontend.scala 304:34]
  assign fq_io_enq_bits_btb_entry = s2_btb_taken ? s2_btb_resp_bits_entry : _GEN_118; // @[Frontend.scala 164:22 Frontend.scala 306:34]
  assign fq_io_enq_bits_btb_bht_history = s2_btb_resp_bits_bht_history; // @[Frontend.scala 164:22]
  assign fq_io_enq_bits_pc = s2_pc; // @[Frontend.scala 158:21]
  assign fq_io_enq_bits_data = icache_io_resp_bits_data; // @[Frontend.scala 161:23]
  assign fq_io_enq_bits_mask = _T_279[1:0]; // @[Frontend.scala 162:23]
  assign fq_io_enq_bits_xcpt_pf_inst = s2_tlb_resp_pf_inst; // @[Frontend.scala 166:23]
  assign fq_io_enq_bits_xcpt_ae_inst = _T_285 | s2_tlb_resp_ae_inst; // @[Frontend.scala 166:23 Frontend.scala 167:87]
  assign fq_io_enq_bits_replay = _T_793 | _GEN_38; // @[Frontend.scala 163:25 Frontend.scala 231:31 Frontend.scala 231:31]
  assign fq_io_deq_ready = io_cpu_resp_ready; // @[Frontend.scala 316:15]
  assign tlb_clock = gated_clock;
  assign tlb_reset = reset;
  assign tlb_io_req_valid = s1_valid & ~s2_replay; // @[Frontend.scala 140:20]
  assign tlb_io_req_bits_vaddr = s1_pc; // @[Frontend.scala 141:25]
  assign tlb_io_sfence_valid = io_cpu_sfence_valid; // @[Frontend.scala 144:17]
  assign tlb_io_sfence_bits_rs1 = io_cpu_sfence_bits_rs1; // @[Frontend.scala 144:17]
  assign tlb_io_sfence_bits_rs2 = io_cpu_sfence_bits_rs2; // @[Frontend.scala 144:17]
  assign tlb_io_sfence_bits_addr = io_cpu_sfence_bits_addr; // @[Frontend.scala 144:17]
  assign tlb_io_ptw_req_ready = io_ptw_req_ready; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_resp_valid = io_ptw_resp_valid; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_resp_bits_ae = io_ptw_resp_bits_ae; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_resp_bits_pte_ppn = io_ptw_resp_bits_pte_ppn; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_resp_bits_pte_d = io_ptw_resp_bits_pte_d; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_resp_bits_pte_a = io_ptw_resp_bits_pte_a; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_resp_bits_pte_g = io_ptw_resp_bits_pte_g; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_resp_bits_pte_u = io_ptw_resp_bits_pte_u; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_resp_bits_pte_x = io_ptw_resp_bits_pte_x; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_resp_bits_pte_w = io_ptw_resp_bits_pte_w; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_resp_bits_pte_r = io_ptw_resp_bits_pte_r; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_resp_bits_pte_v = io_ptw_resp_bits_pte_v; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_resp_bits_level = io_ptw_resp_bits_level; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_resp_bits_homogeneous = io_ptw_resp_bits_homogeneous; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_ptbr_mode = io_ptw_ptbr_mode; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_status_prv = io_ptw_status_prv; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_0_addr = io_ptw_pmp_0_addr; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_0_mask = io_ptw_pmp_0_mask; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_1_addr = io_ptw_pmp_1_addr; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_1_mask = io_ptw_pmp_1_mask; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_2_addr = io_ptw_pmp_2_addr; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_2_mask = io_ptw_pmp_2_mask; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_3_addr = io_ptw_pmp_3_addr; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_3_mask = io_ptw_pmp_3_mask; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_4_addr = io_ptw_pmp_4_addr; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_4_mask = io_ptw_pmp_4_mask; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_5_addr = io_ptw_pmp_5_addr; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_5_mask = io_ptw_pmp_5_mask; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_6_addr = io_ptw_pmp_6_addr; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_6_mask = io_ptw_pmp_6_mask; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_7_addr = io_ptw_pmp_7_addr; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_pmp_7_mask = io_ptw_pmp_7_mask; // @[Frontend.scala 139:10]
  assign tlb_io_ptw_vpoffset_bits_value = io_ptw_vpoffset_bits_value; // @[Frontend.scala 139:10]
  assign tlb_io_kill = ~s2_valid; // @[Frontend.scala 145:15]
  assign btb_clock = gated_clock;
  assign btb_reset = reset;
  assign btb_io_req_bits_addr = s1_pc[38:0]; // @[Frontend.scala 173:26]
  assign btb_io_btb_update_valid = io_cpu_btb_update_valid ? io_cpu_btb_update_valid : _T_303; // @[Frontend.scala 174:23 Frontend.scala 285:31]
  assign btb_io_btb_update_bits_prediction_entry = io_cpu_btb_update_valid ? io_cpu_btb_update_bits_prediction_entry : 5'h1c; // @[Frontend.scala 174:23 Frontend.scala 286:47]
  assign btb_io_btb_update_bits_pc = _GEN_36[38:0]; // @[Frontend.scala 174:23 Frontend.scala 290:33]
  assign btb_io_btb_update_bits_isValid = ~io_cpu_btb_update_valid | io_cpu_btb_update_bits_isValid; // @[Frontend.scala 174:23 Frontend.scala 287:38]
  assign btb_io_btb_update_bits_br_pc = _GEN_35[38:0]; // @[Frontend.scala 174:23 Frontend.scala 289:36]
  assign btb_io_btb_update_bits_cfiType = io_cpu_btb_update_valid ? io_cpu_btb_update_bits_cfiType : btb_io_ras_update_bits_cfiType; // @[Frontend.scala 174:23 Frontend.scala 288:38]
  assign btb_io_bht_update_valid = io_cpu_bht_update_valid; // @[Frontend.scala 175:23 Frontend.scala 190:50]
  assign btb_io_bht_update_bits_prediction_history = io_cpu_bht_update_bits_prediction_history; // @[Frontend.scala 175:23]
  assign btb_io_bht_update_bits_pc = io_cpu_bht_update_bits_pc; // @[Frontend.scala 175:23]
  assign btb_io_bht_update_bits_branch = io_cpu_bht_update_bits_branch; // @[Frontend.scala 175:23]
  assign btb_io_bht_update_bits_taken = io_cpu_bht_update_bits_taken; // @[Frontend.scala 175:23]
  assign btb_io_bht_update_bits_mispredict = io_cpu_bht_update_bits_mispredict; // @[Frontend.scala 175:23]
  assign btb_io_bht_advance_valid = taken_idx ? _GEN_82 : _GEN_46; // @[Frontend.scala 177:30 Frontend.scala 261:36 Frontend.scala 261:36]
  assign btb_io_bht_advance_bits_bht_value = s2_btb_resp_bits_bht_value; // @[Frontend.scala 262:35 Frontend.scala 262:35]
  assign btb_io_ras_update_valid = taken_idx ? _T_803 : _T_536; // @[Frontend.scala 176:29 Frontend.scala 239:33 Frontend.scala 239:33]
  assign btb_io_ras_update_bits_cfiType = taken_idx ? _T_811 : _T_544; // @[Frontend.scala 240:40 Frontend.scala 240:40]
  assign btb_io_ras_update_bits_returnAddr = _T_308[38:0]; // @[Frontend.scala 293:39]
  assign btb_io_flush = _T_793 | _T_526; // @[Frontend.scala 171:18 Frontend.scala 189:54 Frontend.scala 230:22 Frontend.scala 230:22]
  assign Frontend_cov_read_addr = Frontend_state;
  assign Frontend_cov_read_data = Frontend_cov[Frontend_cov_read_addr]; // @[Coverage map for Frontend]
  assign Frontend_cov_write_data = 1'h1;
  assign Frontend_cov_write_addr = Frontend_state;
  assign Frontend_cov_write_mask = 1'h1;
  assign Frontend_cov_write_en = 1'h1;
  assign s2_btb_resp_bits_bht_value_shl = s2_btb_resp_bits_bht_value;
  assign s2_btb_resp_bits_bht_value_pad = {5'h0,s2_btb_resp_bits_bht_value_shl};
  assign s2_btb_resp_bits_taken_shl = {s2_btb_resp_bits_taken, 1'h0};
  assign s2_btb_resp_bits_taken_pad = {4'h0,s2_btb_resp_bits_taken_shl};
  assign _T_249_shl = {_T_249, 2'h0};
  assign _T_249_pad = {3'h0,_T_249_shl};
  assign s2_partial_insn_valid_shl = {s2_partial_insn_valid, 3'h0};
  assign s2_partial_insn_valid_pad = {2'h0,s2_partial_insn_valid_shl};
  assign s2_btb_resp_valid_shl = {s2_btb_resp_valid, 4'h0};
  assign s2_btb_resp_valid_pad = {1'h0,s2_btb_resp_valid_shl};
  assign s2_valid_shl = {s2_valid, 5'h0};
  assign s2_valid_pad = s2_valid_shl;
  assign Frontend_xor4 = s2_btb_resp_bits_taken_pad ^ _T_249_pad;
  assign Frontend_xor1 = s2_btb_resp_bits_bht_value_pad ^ Frontend_xor4;
  assign Frontend_xor6 = s2_btb_resp_valid_pad ^ s2_valid_pad;
  assign Frontend_xor2 = s2_partial_insn_valid_pad ^ Frontend_xor6;
  assign Frontend_xor0 = Frontend_xor1 ^ Frontend_xor2;
  assign icache_sum = Frontend_covSum + icache_io_covSum;
  assign fq_sum = icache_sum + fq_io_covSum;
  assign tlb_sum = fq_sum + tlb_io_covSum;
  assign btb_sum = tlb_sum + btb_io_covSum;
  assign io_covSum = btb_sum;
  assign stopEn0 = ~_T_219;
  assign stopEn1 = ~_T_860;
  assign icache_metaAssert_wire = icache_metaAssert;
  assign fq_metaAssert_wire = fq_metaAssert;
  assign tlb_metaAssert_wire = tlb_metaAssert;
  assign btb_metaAssert_wire = btb_metaAssert;
  assign Frontend_or4 = stopEn1 | icache_metaAssert_wire;
  assign Frontend_or1 = stopEn0 | Frontend_or4;
  assign Frontend_or6 = tlb_metaAssert_wire | btb_metaAssert_wire;
  assign Frontend_or2 = fq_metaAssert_wire | Frontend_or6;
  assign Frontend_or0 = Frontend_or1 | Frontend_or2;
  assign metaAssert = Frontend_or0;
  assign icache_metaReset = metaReset | icache_halt;
  assign fq_metaReset = metaReset | fq_halt;
  assign tlb_metaReset = metaReset | tlb_halt;
  assign btb_metaReset = metaReset | btb_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s1_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  s1_pc = _RAND_1[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  s1_speculative = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  s2_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{`RANDOM}};
  s2_pc = _RAND_4[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  s2_btb_resp_valid = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  s2_btb_resp_bits_taken = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  s2_btb_resp_bits_bridx = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  s2_btb_resp_bits_entry = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  s2_btb_resp_bits_bht_history = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  s2_btb_resp_bits_bht_value = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  s2_tlb_resp_miss = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  s2_tlb_resp_pf_inst = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  s2_tlb_resp_ae_inst = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  s2_tlb_resp_cacheable = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  s2_speculative = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  s2_partial_insn_valid = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  s2_partial_insn = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  wrong_path = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_249 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_268 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  Frontend_state = _RAND_21[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    Frontend_cov[initvar] = _RAND_22[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  Frontend_covSum = _RAND_23[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge gated_clock) begin
    if (metaReset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= io_cpu_req_valid | ~fq_io_mask[2];
    end
    if (metaReset) begin
      s1_pc <= 40'h0;
    end else begin
      s1_pc <= io_cpu_npc;
    end
    if (metaReset) begin
      s1_speculative <= 1'h0;
    end else if (io_cpu_req_valid) begin
      s1_speculative <= io_cpu_req_bits_speculative;
    end else if (s2_replay) begin
      s1_speculative <= s2_speculative;
    end else begin
      s1_speculative <= s0_speculative;
    end
    if (metaReset) begin
      s2_valid <= 1'h0;
    end else if (reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= _GEN_0;
    end
    if (metaReset) begin
      s2_pc <= 40'h0;
    end else if (reset) begin
      s2_pc <= {{8'd0}, ~_T_229};
    end else if (~s2_replay) begin
      s2_pc <= s1_pc;
    end
    if (metaReset) begin
      s2_btb_resp_valid <= 1'h0;
    end else if (~s2_replay) begin
      s2_btb_resp_valid <= btb_io_resp_valid;
    end
    if (metaReset) begin
      s2_btb_resp_bits_taken <= 1'h0;
    end else if (~s2_replay) begin
      s2_btb_resp_bits_taken <= btb_io_resp_bits_taken;
    end
    if (metaReset) begin
      s2_btb_resp_bits_bridx <= 1'h0;
    end else if (~s2_replay) begin
      s2_btb_resp_bits_bridx <= btb_io_resp_bits_bridx;
    end
    if (metaReset) begin
      s2_btb_resp_bits_entry <= 5'h0;
    end else if (~s2_replay) begin
      s2_btb_resp_bits_entry <= btb_io_resp_bits_entry;
    end
    if (metaReset) begin
      s2_btb_resp_bits_bht_history <= 8'h0;
    end else if (~s2_replay) begin
      s2_btb_resp_bits_bht_history <= btb_io_resp_bits_bht_history;
    end
    if (metaReset) begin
      s2_btb_resp_bits_bht_value <= 1'h0;
    end else if (~s2_replay) begin
      s2_btb_resp_bits_bht_value <= btb_io_resp_bits_bht_value;
    end
    if (metaReset) begin
      s2_tlb_resp_miss <= 1'h0;
    end else if (~s2_replay) begin
      s2_tlb_resp_miss <= tlb_io_resp_miss;
    end
    if (metaReset) begin
      s2_tlb_resp_pf_inst <= 1'h0;
    end else if (~s2_replay) begin
      s2_tlb_resp_pf_inst <= tlb_io_resp_pf_inst;
    end
    if (metaReset) begin
      s2_tlb_resp_ae_inst <= 1'h0;
    end else if (~s2_replay) begin
      s2_tlb_resp_ae_inst <= tlb_io_resp_ae_inst;
    end
    if (metaReset) begin
      s2_tlb_resp_cacheable <= 1'h0;
    end else if (~s2_replay) begin
      s2_tlb_resp_cacheable <= tlb_io_resp_cacheable;
    end
    if (metaReset) begin
      s2_speculative <= 1'h0;
    end else if (reset) begin
      s2_speculative <= 1'h0;
    end else if (~s2_replay) begin
      s2_speculative <= s1_speculative;
    end
    if (metaReset) begin
      s2_partial_insn_valid <= 1'h0;
    end else if (reset) begin
      s2_partial_insn_valid <= 1'h0;
    end else if (s2_redirect) begin
      s2_partial_insn_valid <= 1'h0;
    end else if (_T_853) begin
      s2_partial_insn_valid <= 1'h0;
    end else if (_T_243) begin
      s2_partial_insn_valid <= _T_849;
    end
    if (metaReset) begin
      s2_partial_insn <= 16'h0;
    end else if (_T_243) begin
      if (_T_849) begin
        s2_partial_insn <= _T_850;
      end
    end
    if (metaReset) begin
      wrong_path <= 1'h0;
    end else if (io_cpu_req_valid) begin
      wrong_path <= 1'h0;
    end else if (taken_idx) begin
      if (~s2_btb_taken) begin
        wrong_path <= _GEN_76;
      end else begin
        wrong_path <= _GEN_75;
      end
    end else begin
      wrong_path <= _GEN_75;
    end
    if (metaReset) begin
      _T_249 <= 1'h0;
    end else begin
      _T_249 <= reset | _T_247;
    end
    if (metaReset) begin
      _T_268 <= 1'h0;
    end else begin
      _T_268 <= s1_valid;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_219) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Frontend.scala:86 assert(!(io.cpu.req.valid || io.cpu.sfence.valid || io.cpu.flush_icache || io.cpu.bht_update.valid || io.cpu.btb_update.valid) || io.cpu.might_request)\n"); // @[Frontend.scala 86:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_219) begin
          $fatal; // @[Frontend.scala 86:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_860) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Frontend.scala:311 assert(!s2_partial_insn_valid || fq.io.enq.bits.mask(0))\n"); // @[Frontend.scala 311:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_860) begin
          $fatal; // @[Frontend.scala 311:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    Frontend_state <= Frontend_xor0;
    if (!(Frontend_cov_read_data)) begin
      Frontend_covSum <= Frontend_covSum + 1'h1;
    end
  end
  always @(posedge gated_clock) begin
    if(Frontend_cov_write_en & Frontend_cov_write_mask) begin
      Frontend_cov[Frontend_cov_write_addr] <= Frontend_cov_write_data; // @[Coverage map for Frontend]
    end
  end
endmodule
module TLBuffer_22(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [3:0]  auto_in_a_bits_size,
  input  [1:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_a_bits_corrupt,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [2:0]  auto_in_b_bits_opcode,
  output [1:0]  auto_in_b_bits_param,
  output [3:0]  auto_in_b_bits_size,
  output [1:0]  auto_in_b_bits_source,
  output [31:0] auto_in_b_bits_address,
  output [7:0]  auto_in_b_bits_mask,
  output        auto_in_b_bits_corrupt,
  output        auto_in_c_ready,
  input         auto_in_c_valid,
  input  [2:0]  auto_in_c_bits_opcode,
  input  [2:0]  auto_in_c_bits_param,
  input  [3:0]  auto_in_c_bits_size,
  input  [1:0]  auto_in_c_bits_source,
  input  [31:0] auto_in_c_bits_address,
  input  [63:0] auto_in_c_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [1:0]  auto_in_d_bits_param,
  output [3:0]  auto_in_d_bits_size,
  output [1:0]  auto_in_d_bits_source,
  output [1:0]  auto_in_d_bits_sink,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  output        auto_in_e_ready,
  input         auto_in_e_valid,
  input  [1:0]  auto_in_e_bits_sink,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [3:0]  auto_out_a_bits_size,
  output [1:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_a_bits_corrupt,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [2:0]  auto_out_b_bits_opcode,
  input  [1:0]  auto_out_b_bits_param,
  input  [3:0]  auto_out_b_bits_size,
  input  [1:0]  auto_out_b_bits_source,
  input  [31:0] auto_out_b_bits_address,
  input  [7:0]  auto_out_b_bits_mask,
  input         auto_out_b_bits_corrupt,
  input         auto_out_c_ready,
  output        auto_out_c_valid,
  output [2:0]  auto_out_c_bits_opcode,
  output [2:0]  auto_out_c_bits_param,
  output [3:0]  auto_out_c_bits_size,
  output [1:0]  auto_out_c_bits_source,
  output [31:0] auto_out_c_bits_address,
  output [63:0] auto_out_c_bits_data,
  output        auto_out_c_bits_corrupt,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_param,
  input  [3:0]  auto_out_d_bits_size,
  input  [1:0]  auto_out_d_bits_source,
  input  [1:0]  auto_out_d_bits_sink,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  input         auto_out_e_ready,
  output        auto_out_e_valid,
  output [1:0]  auto_out_e_bits_sink,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         TLMonitor_halt,
  input         Queue_4_halt,
  input         Queue_2_halt,
  input         Queue_1_halt,
  input         Queue_3_halt,
  input         Queue_halt
);
  wire  TLMonitor_clock; // @[Nodes.scala 25:25]
  wire  TLMonitor_reset; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_a_ready; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_a_valid; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_a_bits_opcode; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_a_bits_param; // @[Nodes.scala 25:25]
  wire [3:0] TLMonitor_io_in_a_bits_size; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_a_bits_source; // @[Nodes.scala 25:25]
  wire [31:0] TLMonitor_io_in_a_bits_address; // @[Nodes.scala 25:25]
  wire [7:0] TLMonitor_io_in_a_bits_mask; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_a_bits_corrupt; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_b_ready; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_b_valid; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_b_bits_opcode; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_b_bits_param; // @[Nodes.scala 25:25]
  wire [3:0] TLMonitor_io_in_b_bits_size; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_b_bits_source; // @[Nodes.scala 25:25]
  wire [31:0] TLMonitor_io_in_b_bits_address; // @[Nodes.scala 25:25]
  wire [7:0] TLMonitor_io_in_b_bits_mask; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_b_bits_corrupt; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_c_ready; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_c_valid; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_c_bits_opcode; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_c_bits_param; // @[Nodes.scala 25:25]
  wire [3:0] TLMonitor_io_in_c_bits_size; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_c_bits_source; // @[Nodes.scala 25:25]
  wire [31:0] TLMonitor_io_in_c_bits_address; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_d_ready; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_d_valid; // @[Nodes.scala 25:25]
  wire [2:0] TLMonitor_io_in_d_bits_opcode; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_d_bits_param; // @[Nodes.scala 25:25]
  wire [3:0] TLMonitor_io_in_d_bits_size; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_d_bits_source; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_d_bits_sink; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_d_bits_denied; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_d_bits_corrupt; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_e_ready; // @[Nodes.scala 25:25]
  wire  TLMonitor_io_in_e_valid; // @[Nodes.scala 25:25]
  wire [1:0] TLMonitor_io_in_e_bits_sink; // @[Nodes.scala 25:25]
  wire [29:0] TLMonitor_io_covSum; // @[Nodes.scala 25:25]
  wire  TLMonitor_metaAssert; // @[Nodes.scala 25:25]
  wire  TLMonitor_metaReset; // @[Nodes.scala 25:25]
  wire  Queue_clock; // @[Decoupled.scala 293:21]
  wire  Queue_reset; // @[Decoupled.scala 293:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 293:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 293:21]
  wire [2:0] Queue_io_enq_bits_opcode; // @[Decoupled.scala 293:21]
  wire [2:0] Queue_io_enq_bits_param; // @[Decoupled.scala 293:21]
  wire [3:0] Queue_io_enq_bits_size; // @[Decoupled.scala 293:21]
  wire [1:0] Queue_io_enq_bits_source; // @[Decoupled.scala 293:21]
  wire [31:0] Queue_io_enq_bits_address; // @[Decoupled.scala 293:21]
  wire [7:0] Queue_io_enq_bits_mask; // @[Decoupled.scala 293:21]
  wire [63:0] Queue_io_enq_bits_data; // @[Decoupled.scala 293:21]
  wire  Queue_io_enq_bits_corrupt; // @[Decoupled.scala 293:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 293:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 293:21]
  wire [2:0] Queue_io_deq_bits_opcode; // @[Decoupled.scala 293:21]
  wire [2:0] Queue_io_deq_bits_param; // @[Decoupled.scala 293:21]
  wire [3:0] Queue_io_deq_bits_size; // @[Decoupled.scala 293:21]
  wire [1:0] Queue_io_deq_bits_source; // @[Decoupled.scala 293:21]
  wire [31:0] Queue_io_deq_bits_address; // @[Decoupled.scala 293:21]
  wire [7:0] Queue_io_deq_bits_mask; // @[Decoupled.scala 293:21]
  wire [63:0] Queue_io_deq_bits_data; // @[Decoupled.scala 293:21]
  wire  Queue_io_deq_bits_corrupt; // @[Decoupled.scala 293:21]
  wire [29:0] Queue_io_covSum; // @[Decoupled.scala 293:21]
  wire  Queue_metaAssert; // @[Decoupled.scala 293:21]
  wire  Queue_metaReset; // @[Decoupled.scala 293:21]
  wire  Queue_1_clock; // @[Decoupled.scala 293:21]
  wire  Queue_1_reset; // @[Decoupled.scala 293:21]
  wire  Queue_1_io_enq_ready; // @[Decoupled.scala 293:21]
  wire  Queue_1_io_enq_valid; // @[Decoupled.scala 293:21]
  wire [2:0] Queue_1_io_enq_bits_opcode; // @[Decoupled.scala 293:21]
  wire [1:0] Queue_1_io_enq_bits_param; // @[Decoupled.scala 293:21]
  wire [3:0] Queue_1_io_enq_bits_size; // @[Decoupled.scala 293:21]
  wire [1:0] Queue_1_io_enq_bits_source; // @[Decoupled.scala 293:21]
  wire [1:0] Queue_1_io_enq_bits_sink; // @[Decoupled.scala 293:21]
  wire  Queue_1_io_enq_bits_denied; // @[Decoupled.scala 293:21]
  wire [63:0] Queue_1_io_enq_bits_data; // @[Decoupled.scala 293:21]
  wire  Queue_1_io_enq_bits_corrupt; // @[Decoupled.scala 293:21]
  wire  Queue_1_io_deq_ready; // @[Decoupled.scala 293:21]
  wire  Queue_1_io_deq_valid; // @[Decoupled.scala 293:21]
  wire [2:0] Queue_1_io_deq_bits_opcode; // @[Decoupled.scala 293:21]
  wire [1:0] Queue_1_io_deq_bits_param; // @[Decoupled.scala 293:21]
  wire [3:0] Queue_1_io_deq_bits_size; // @[Decoupled.scala 293:21]
  wire [1:0] Queue_1_io_deq_bits_source; // @[Decoupled.scala 293:21]
  wire [1:0] Queue_1_io_deq_bits_sink; // @[Decoupled.scala 293:21]
  wire  Queue_1_io_deq_bits_denied; // @[Decoupled.scala 293:21]
  wire [63:0] Queue_1_io_deq_bits_data; // @[Decoupled.scala 293:21]
  wire  Queue_1_io_deq_bits_corrupt; // @[Decoupled.scala 293:21]
  wire [29:0] Queue_1_io_covSum; // @[Decoupled.scala 293:21]
  wire  Queue_1_metaAssert; // @[Decoupled.scala 293:21]
  wire  Queue_1_metaReset; // @[Decoupled.scala 293:21]
  wire  Queue_2_clock; // @[Decoupled.scala 293:21]
  wire  Queue_2_reset; // @[Decoupled.scala 293:21]
  wire  Queue_2_io_enq_ready; // @[Decoupled.scala 293:21]
  wire  Queue_2_io_enq_valid; // @[Decoupled.scala 293:21]
  wire [2:0] Queue_2_io_enq_bits_opcode; // @[Decoupled.scala 293:21]
  wire [1:0] Queue_2_io_enq_bits_param; // @[Decoupled.scala 293:21]
  wire [3:0] Queue_2_io_enq_bits_size; // @[Decoupled.scala 293:21]
  wire [1:0] Queue_2_io_enq_bits_source; // @[Decoupled.scala 293:21]
  wire [31:0] Queue_2_io_enq_bits_address; // @[Decoupled.scala 293:21]
  wire [7:0] Queue_2_io_enq_bits_mask; // @[Decoupled.scala 293:21]
  wire  Queue_2_io_enq_bits_corrupt; // @[Decoupled.scala 293:21]
  wire  Queue_2_io_deq_ready; // @[Decoupled.scala 293:21]
  wire  Queue_2_io_deq_valid; // @[Decoupled.scala 293:21]
  wire [2:0] Queue_2_io_deq_bits_opcode; // @[Decoupled.scala 293:21]
  wire [1:0] Queue_2_io_deq_bits_param; // @[Decoupled.scala 293:21]
  wire [3:0] Queue_2_io_deq_bits_size; // @[Decoupled.scala 293:21]
  wire [1:0] Queue_2_io_deq_bits_source; // @[Decoupled.scala 293:21]
  wire [31:0] Queue_2_io_deq_bits_address; // @[Decoupled.scala 293:21]
  wire [7:0] Queue_2_io_deq_bits_mask; // @[Decoupled.scala 293:21]
  wire  Queue_2_io_deq_bits_corrupt; // @[Decoupled.scala 293:21]
  wire [29:0] Queue_2_io_covSum; // @[Decoupled.scala 293:21]
  wire  Queue_2_metaAssert; // @[Decoupled.scala 293:21]
  wire  Queue_2_metaReset; // @[Decoupled.scala 293:21]
  wire  Queue_3_clock; // @[Decoupled.scala 293:21]
  wire  Queue_3_reset; // @[Decoupled.scala 293:21]
  wire  Queue_3_io_enq_ready; // @[Decoupled.scala 293:21]
  wire  Queue_3_io_enq_valid; // @[Decoupled.scala 293:21]
  wire [2:0] Queue_3_io_enq_bits_opcode; // @[Decoupled.scala 293:21]
  wire [2:0] Queue_3_io_enq_bits_param; // @[Decoupled.scala 293:21]
  wire [3:0] Queue_3_io_enq_bits_size; // @[Decoupled.scala 293:21]
  wire [1:0] Queue_3_io_enq_bits_source; // @[Decoupled.scala 293:21]
  wire [31:0] Queue_3_io_enq_bits_address; // @[Decoupled.scala 293:21]
  wire [63:0] Queue_3_io_enq_bits_data; // @[Decoupled.scala 293:21]
  wire  Queue_3_io_deq_ready; // @[Decoupled.scala 293:21]
  wire  Queue_3_io_deq_valid; // @[Decoupled.scala 293:21]
  wire [2:0] Queue_3_io_deq_bits_opcode; // @[Decoupled.scala 293:21]
  wire [2:0] Queue_3_io_deq_bits_param; // @[Decoupled.scala 293:21]
  wire [3:0] Queue_3_io_deq_bits_size; // @[Decoupled.scala 293:21]
  wire [1:0] Queue_3_io_deq_bits_source; // @[Decoupled.scala 293:21]
  wire [31:0] Queue_3_io_deq_bits_address; // @[Decoupled.scala 293:21]
  wire [63:0] Queue_3_io_deq_bits_data; // @[Decoupled.scala 293:21]
  wire  Queue_3_io_deq_bits_corrupt; // @[Decoupled.scala 293:21]
  wire [29:0] Queue_3_io_covSum; // @[Decoupled.scala 293:21]
  wire  Queue_3_metaAssert; // @[Decoupled.scala 293:21]
  wire  Queue_3_metaReset; // @[Decoupled.scala 293:21]
  wire  Queue_4_clock; // @[Decoupled.scala 293:21]
  wire  Queue_4_reset; // @[Decoupled.scala 293:21]
  wire  Queue_4_io_enq_ready; // @[Decoupled.scala 293:21]
  wire  Queue_4_io_enq_valid; // @[Decoupled.scala 293:21]
  wire [1:0] Queue_4_io_enq_bits_sink; // @[Decoupled.scala 293:21]
  wire  Queue_4_io_deq_ready; // @[Decoupled.scala 293:21]
  wire  Queue_4_io_deq_valid; // @[Decoupled.scala 293:21]
  wire [1:0] Queue_4_io_deq_bits_sink; // @[Decoupled.scala 293:21]
  wire [29:0] Queue_4_io_covSum; // @[Decoupled.scala 293:21]
  wire  Queue_4_metaAssert; // @[Decoupled.scala 293:21]
  wire  Queue_4_metaReset; // @[Decoupled.scala 293:21]
  wire [29:0] TLBuffer_22_covSum;
  wire [29:0] TLMonitor_sum;
  wire [29:0] Queue_4_sum;
  wire [29:0] Queue_2_sum;
  wire [29:0] Queue_1_sum;
  wire [29:0] Queue_3_sum;
  wire [29:0] Queue_sum;
  wire  TLMonitor_metaAssert_wire;
  wire  Queue_metaAssert_wire;
  wire  Queue_1_metaAssert_wire;
  wire  Queue_4_metaAssert_wire;
  wire  Queue_3_metaAssert_wire;
  wire  Queue_2_metaAssert_wire;
  wire  TLBuffer_22_or4;
  wire  TLBuffer_22_or1;
  wire  TLBuffer_22_or6;
  wire  TLBuffer_22_or2;
  wire  TLBuffer_22_or0;
  reg  TLBuffer_22_metaAssert;
  reg [31:0] _RAND_0;
  TLMonitor_66 TLMonitor ( // @[Nodes.scala 25:25]
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_io_in_a_bits_corrupt),
    .io_in_b_ready(TLMonitor_io_in_b_ready),
    .io_in_b_valid(TLMonitor_io_in_b_valid),
    .io_in_b_bits_opcode(TLMonitor_io_in_b_bits_opcode),
    .io_in_b_bits_param(TLMonitor_io_in_b_bits_param),
    .io_in_b_bits_size(TLMonitor_io_in_b_bits_size),
    .io_in_b_bits_source(TLMonitor_io_in_b_bits_source),
    .io_in_b_bits_address(TLMonitor_io_in_b_bits_address),
    .io_in_b_bits_mask(TLMonitor_io_in_b_bits_mask),
    .io_in_b_bits_corrupt(TLMonitor_io_in_b_bits_corrupt),
    .io_in_c_ready(TLMonitor_io_in_c_ready),
    .io_in_c_valid(TLMonitor_io_in_c_valid),
    .io_in_c_bits_opcode(TLMonitor_io_in_c_bits_opcode),
    .io_in_c_bits_param(TLMonitor_io_in_c_bits_param),
    .io_in_c_bits_size(TLMonitor_io_in_c_bits_size),
    .io_in_c_bits_source(TLMonitor_io_in_c_bits_source),
    .io_in_c_bits_address(TLMonitor_io_in_c_bits_address),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt),
    .io_in_e_ready(TLMonitor_io_in_e_ready),
    .io_in_e_valid(TLMonitor_io_in_e_valid),
    .io_in_e_bits_sink(TLMonitor_io_in_e_bits_sink),
    .io_covSum(TLMonitor_io_covSum),
    .metaAssert(TLMonitor_metaAssert),
    .metaReset(TLMonitor_metaReset)
  );
  Queue_108 Queue ( // @[Decoupled.scala 293:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_opcode(Queue_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_io_enq_bits_param),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_enq_bits_source(Queue_io_enq_bits_source),
    .io_enq_bits_address(Queue_io_enq_bits_address),
    .io_enq_bits_mask(Queue_io_enq_bits_mask),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_corrupt(Queue_io_enq_bits_corrupt),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_opcode(Queue_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_io_deq_bits_param),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_source(Queue_io_deq_bits_source),
    .io_deq_bits_address(Queue_io_deq_bits_address),
    .io_deq_bits_mask(Queue_io_deq_bits_mask),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_corrupt(Queue_io_deq_bits_corrupt),
    .io_covSum(Queue_io_covSum),
    .metaAssert(Queue_metaAssert),
    .metaReset(Queue_metaReset)
  );
  Queue_109 Queue_1 ( // @[Decoupled.scala 293:21]
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_opcode(Queue_1_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_1_io_enq_bits_param),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_source(Queue_1_io_enq_bits_source),
    .io_enq_bits_sink(Queue_1_io_enq_bits_sink),
    .io_enq_bits_denied(Queue_1_io_enq_bits_denied),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_corrupt(Queue_1_io_enq_bits_corrupt),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_opcode(Queue_1_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_1_io_deq_bits_param),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_source(Queue_1_io_deq_bits_source),
    .io_deq_bits_sink(Queue_1_io_deq_bits_sink),
    .io_deq_bits_denied(Queue_1_io_deq_bits_denied),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_corrupt(Queue_1_io_deq_bits_corrupt),
    .io_covSum(Queue_1_io_covSum),
    .metaAssert(Queue_1_metaAssert),
    .metaReset(Queue_1_metaReset)
  );
  Queue_110 Queue_2 ( // @[Decoupled.scala 293:21]
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_opcode(Queue_2_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_2_io_enq_bits_param),
    .io_enq_bits_size(Queue_2_io_enq_bits_size),
    .io_enq_bits_source(Queue_2_io_enq_bits_source),
    .io_enq_bits_address(Queue_2_io_enq_bits_address),
    .io_enq_bits_mask(Queue_2_io_enq_bits_mask),
    .io_enq_bits_corrupt(Queue_2_io_enq_bits_corrupt),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_opcode(Queue_2_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_2_io_deq_bits_param),
    .io_deq_bits_size(Queue_2_io_deq_bits_size),
    .io_deq_bits_source(Queue_2_io_deq_bits_source),
    .io_deq_bits_address(Queue_2_io_deq_bits_address),
    .io_deq_bits_mask(Queue_2_io_deq_bits_mask),
    .io_deq_bits_corrupt(Queue_2_io_deq_bits_corrupt),
    .io_covSum(Queue_2_io_covSum),
    .metaAssert(Queue_2_metaAssert),
    .metaReset(Queue_2_metaReset)
  );
  Queue_111 Queue_3 ( // @[Decoupled.scala 293:21]
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits_opcode(Queue_3_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_3_io_enq_bits_param),
    .io_enq_bits_size(Queue_3_io_enq_bits_size),
    .io_enq_bits_source(Queue_3_io_enq_bits_source),
    .io_enq_bits_address(Queue_3_io_enq_bits_address),
    .io_enq_bits_data(Queue_3_io_enq_bits_data),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits_opcode(Queue_3_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_3_io_deq_bits_param),
    .io_deq_bits_size(Queue_3_io_deq_bits_size),
    .io_deq_bits_source(Queue_3_io_deq_bits_source),
    .io_deq_bits_address(Queue_3_io_deq_bits_address),
    .io_deq_bits_data(Queue_3_io_deq_bits_data),
    .io_deq_bits_corrupt(Queue_3_io_deq_bits_corrupt),
    .io_covSum(Queue_3_io_covSum),
    .metaAssert(Queue_3_metaAssert),
    .metaReset(Queue_3_metaReset)
  );
  Queue_112 Queue_4 ( // @[Decoupled.scala 293:21]
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits_sink(Queue_4_io_enq_bits_sink),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits_sink(Queue_4_io_deq_bits_sink),
    .io_covSum(Queue_4_io_covSum),
    .metaAssert(Queue_4_metaAssert),
    .metaReset(Queue_4_metaReset)
  );
  assign auto_in_a_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_in_b_valid = Queue_2_io_deq_valid; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_opcode = Queue_2_io_deq_bits_opcode; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_param = Queue_2_io_deq_bits_param; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_size = Queue_2_io_deq_bits_size; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_source = Queue_2_io_deq_bits_source; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_address = Queue_2_io_deq_bits_address; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_mask = Queue_2_io_deq_bits_mask; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_corrupt = Queue_2_io_deq_bits_corrupt; // @[LazyModule.scala 173:31]
  assign auto_in_c_ready = Queue_3_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_in_d_valid = Queue_1_io_deq_valid; // @[LazyModule.scala 173:31]
  assign auto_in_d_bits_opcode = Queue_1_io_deq_bits_opcode; // @[LazyModule.scala 173:31]
  assign auto_in_d_bits_param = Queue_1_io_deq_bits_param; // @[LazyModule.scala 173:31]
  assign auto_in_d_bits_size = Queue_1_io_deq_bits_size; // @[LazyModule.scala 173:31]
  assign auto_in_d_bits_source = Queue_1_io_deq_bits_source; // @[LazyModule.scala 173:31]
  assign auto_in_d_bits_sink = Queue_1_io_deq_bits_sink; // @[LazyModule.scala 173:31]
  assign auto_in_d_bits_denied = Queue_1_io_deq_bits_denied; // @[LazyModule.scala 173:31]
  assign auto_in_d_bits_data = Queue_1_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_in_d_bits_corrupt = Queue_1_io_deq_bits_corrupt; // @[LazyModule.scala 173:31]
  assign auto_in_e_ready = Queue_4_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_out_a_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_opcode = Queue_io_deq_bits_opcode; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_param = Queue_io_deq_bits_param; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_size = Queue_io_deq_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_source = Queue_io_deq_bits_source; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_address = Queue_io_deq_bits_address; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_mask = Queue_io_deq_bits_mask; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_a_bits_corrupt = Queue_io_deq_bits_corrupt; // @[LazyModule.scala 173:49]
  assign auto_out_b_ready = Queue_2_io_enq_ready; // @[LazyModule.scala 173:49]
  assign auto_out_c_valid = Queue_3_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_c_bits_opcode = Queue_3_io_deq_bits_opcode; // @[LazyModule.scala 173:49]
  assign auto_out_c_bits_param = Queue_3_io_deq_bits_param; // @[LazyModule.scala 173:49]
  assign auto_out_c_bits_size = Queue_3_io_deq_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_c_bits_source = Queue_3_io_deq_bits_source; // @[LazyModule.scala 173:49]
  assign auto_out_c_bits_address = Queue_3_io_deq_bits_address; // @[LazyModule.scala 173:49]
  assign auto_out_c_bits_data = Queue_3_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_c_bits_corrupt = Queue_3_io_deq_bits_corrupt; // @[LazyModule.scala 173:49]
  assign auto_out_d_ready = Queue_1_io_enq_ready; // @[LazyModule.scala 173:49]
  assign auto_out_e_valid = Queue_4_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_e_bits_sink = Queue_4_io_deq_bits_sink; // @[LazyModule.scala 173:49]
  assign TLMonitor_clock = clock;
  assign TLMonitor_reset = reset;
  assign TLMonitor_io_in_a_ready = Queue_io_enq_ready; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_ready = auto_in_b_ready; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_valid = Queue_2_io_deq_valid; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_opcode = Queue_2_io_deq_bits_opcode; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_param = Queue_2_io_deq_bits_param; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_size = Queue_2_io_deq_bits_size; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_source = Queue_2_io_deq_bits_source; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_address = Queue_2_io_deq_bits_address; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_mask = Queue_2_io_deq_bits_mask; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_b_bits_corrupt = Queue_2_io_deq_bits_corrupt; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_ready = Queue_3_io_enq_ready; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_valid = auto_in_c_valid; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_bits_opcode = auto_in_c_bits_opcode; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_bits_param = auto_in_c_bits_param; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_bits_size = auto_in_c_bits_size; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_bits_source = auto_in_c_bits_source; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_c_bits_address = auto_in_c_bits_address; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_valid = Queue_1_io_deq_valid; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_opcode = Queue_1_io_deq_bits_opcode; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_param = Queue_1_io_deq_bits_param; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_size = Queue_1_io_deq_bits_size; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_source = Queue_1_io_deq_bits_source; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_sink = Queue_1_io_deq_bits_sink; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_denied = Queue_1_io_deq_bits_denied; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_d_bits_corrupt = Queue_1_io_deq_bits_corrupt; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_e_ready = Queue_4_io_enq_ready; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_e_valid = auto_in_e_valid; // @[Nodes.scala 26:19]
  assign TLMonitor_io_in_e_bits_sink = auto_in_e_bits_sink; // @[Nodes.scala 26:19]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_a_valid; // @[Decoupled.scala 294:22]
  assign Queue_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Decoupled.scala 295:21]
  assign Queue_io_enq_bits_param = auto_in_a_bits_param; // @[Decoupled.scala 295:21]
  assign Queue_io_enq_bits_size = auto_in_a_bits_size; // @[Decoupled.scala 295:21]
  assign Queue_io_enq_bits_source = auto_in_a_bits_source; // @[Decoupled.scala 295:21]
  assign Queue_io_enq_bits_address = auto_in_a_bits_address; // @[Decoupled.scala 295:21]
  assign Queue_io_enq_bits_mask = auto_in_a_bits_mask; // @[Decoupled.scala 295:21]
  assign Queue_io_enq_bits_data = auto_in_a_bits_data; // @[Decoupled.scala 295:21]
  assign Queue_io_enq_bits_corrupt = auto_in_a_bits_corrupt; // @[Decoupled.scala 295:21]
  assign Queue_io_deq_ready = auto_out_a_ready; // @[Buffer.scala 38:13]
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = auto_out_d_valid; // @[Decoupled.scala 294:22]
  assign Queue_1_io_enq_bits_opcode = auto_out_d_bits_opcode; // @[Decoupled.scala 295:21]
  assign Queue_1_io_enq_bits_param = auto_out_d_bits_param; // @[Decoupled.scala 295:21]
  assign Queue_1_io_enq_bits_size = auto_out_d_bits_size; // @[Decoupled.scala 295:21]
  assign Queue_1_io_enq_bits_source = auto_out_d_bits_source; // @[Decoupled.scala 295:21]
  assign Queue_1_io_enq_bits_sink = auto_out_d_bits_sink; // @[Decoupled.scala 295:21]
  assign Queue_1_io_enq_bits_denied = auto_out_d_bits_denied; // @[Decoupled.scala 295:21]
  assign Queue_1_io_enq_bits_data = auto_out_d_bits_data; // @[Decoupled.scala 295:21]
  assign Queue_1_io_enq_bits_corrupt = auto_out_d_bits_corrupt; // @[Decoupled.scala 295:21]
  assign Queue_1_io_deq_ready = auto_in_d_ready; // @[Buffer.scala 39:13]
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_2_io_enq_valid = auto_out_b_valid; // @[Decoupled.scala 294:22]
  assign Queue_2_io_enq_bits_opcode = auto_out_b_bits_opcode; // @[Decoupled.scala 295:21]
  assign Queue_2_io_enq_bits_param = auto_out_b_bits_param; // @[Decoupled.scala 295:21]
  assign Queue_2_io_enq_bits_size = auto_out_b_bits_size; // @[Decoupled.scala 295:21]
  assign Queue_2_io_enq_bits_source = auto_out_b_bits_source; // @[Decoupled.scala 295:21]
  assign Queue_2_io_enq_bits_address = auto_out_b_bits_address; // @[Decoupled.scala 295:21]
  assign Queue_2_io_enq_bits_mask = auto_out_b_bits_mask; // @[Decoupled.scala 295:21]
  assign Queue_2_io_enq_bits_corrupt = auto_out_b_bits_corrupt; // @[Decoupled.scala 295:21]
  assign Queue_2_io_deq_ready = auto_in_b_ready; // @[Buffer.scala 42:15]
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign Queue_3_io_enq_valid = auto_in_c_valid; // @[Decoupled.scala 294:22]
  assign Queue_3_io_enq_bits_opcode = auto_in_c_bits_opcode; // @[Decoupled.scala 295:21]
  assign Queue_3_io_enq_bits_param = auto_in_c_bits_param; // @[Decoupled.scala 295:21]
  assign Queue_3_io_enq_bits_size = auto_in_c_bits_size; // @[Decoupled.scala 295:21]
  assign Queue_3_io_enq_bits_source = auto_in_c_bits_source; // @[Decoupled.scala 295:21]
  assign Queue_3_io_enq_bits_address = auto_in_c_bits_address; // @[Decoupled.scala 295:21]
  assign Queue_3_io_enq_bits_data = auto_in_c_bits_data; // @[Decoupled.scala 295:21]
  assign Queue_3_io_deq_ready = auto_out_c_ready; // @[Buffer.scala 43:15]
  assign Queue_4_clock = clock;
  assign Queue_4_reset = reset;
  assign Queue_4_io_enq_valid = auto_in_e_valid; // @[Decoupled.scala 294:22]
  assign Queue_4_io_enq_bits_sink = auto_in_e_bits_sink; // @[Decoupled.scala 295:21]
  assign Queue_4_io_deq_ready = auto_out_e_ready; // @[Buffer.scala 44:15]
  assign TLBuffer_22_covSum = 30'h0;
  assign TLMonitor_sum = TLBuffer_22_covSum + TLMonitor_io_covSum;
  assign Queue_4_sum = TLMonitor_sum + Queue_4_io_covSum;
  assign Queue_2_sum = Queue_4_sum + Queue_2_io_covSum;
  assign Queue_1_sum = Queue_2_sum + Queue_1_io_covSum;
  assign Queue_3_sum = Queue_1_sum + Queue_3_io_covSum;
  assign Queue_sum = Queue_3_sum + Queue_io_covSum;
  assign io_covSum = Queue_sum;
  assign TLMonitor_metaAssert_wire = TLMonitor_metaAssert;
  assign Queue_2_metaAssert_wire = Queue_2_metaAssert;
  assign Queue_4_metaAssert_wire = Queue_4_metaAssert;
  assign Queue_1_metaAssert_wire = Queue_1_metaAssert;
  assign Queue_metaAssert_wire = Queue_metaAssert;
  assign Queue_3_metaAssert_wire = Queue_3_metaAssert;
  assign TLBuffer_22_or4 = Queue_4_metaAssert_wire | TLMonitor_metaAssert_wire;
  assign TLBuffer_22_or1 = Queue_2_metaAssert_wire | TLBuffer_22_or4;
  assign TLBuffer_22_or6 = Queue_metaAssert_wire | Queue_3_metaAssert_wire;
  assign TLBuffer_22_or2 = Queue_1_metaAssert_wire | TLBuffer_22_or6;
  assign TLBuffer_22_or0 = TLBuffer_22_or1 | TLBuffer_22_or2;
  assign metaAssert = TLBuffer_22_metaAssert;
  assign TLMonitor_metaReset = metaReset | TLMonitor_halt;
  assign Queue_4_metaReset = metaReset | Queue_4_halt;
  assign Queue_2_metaReset = metaReset | Queue_2_halt;
  assign Queue_1_metaReset = metaReset | Queue_1_halt;
  assign Queue_3_metaReset = metaReset | Queue_3_halt;
  assign Queue_metaReset = metaReset | Queue_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  TLBuffer_22_metaAssert = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      TLBuffer_22_metaAssert <= 1'h0;
    end else begin
      TLBuffer_22_metaAssert <= TLBuffer_22_metaAssert | TLBuffer_22_or0;
    end
  end
endmodule
module IntSyncCrossingSink(
  input         clock,
  input         auto_in_sync_0,
  output        auto_out_0,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         SynchronizerShiftReg_w1_d3_halt
);
  wire  SynchronizerShiftReg_w1_d3_clock; // @[ShiftReg.scala 47:23]
  wire  SynchronizerShiftReg_w1_d3_io_d; // @[ShiftReg.scala 47:23]
  wire  SynchronizerShiftReg_w1_d3_io_q; // @[ShiftReg.scala 47:23]
  wire [29:0] SynchronizerShiftReg_w1_d3_io_covSum; // @[ShiftReg.scala 47:23]
  wire  SynchronizerShiftReg_w1_d3_metaAssert; // @[ShiftReg.scala 47:23]
  wire  SynchronizerShiftReg_w1_d3_metaReset; // @[ShiftReg.scala 47:23]
  wire [29:0] IntSyncCrossingSink_covSum;
  wire [29:0] SynchronizerShiftReg_w1_d3_sum;
  wire  SynchronizerShiftReg_w1_d3_metaAssert_wire;
  SynchronizerShiftReg_w1_d3 SynchronizerShiftReg_w1_d3 ( // @[ShiftReg.scala 47:23]
    .clock(SynchronizerShiftReg_w1_d3_clock),
    .io_d(SynchronizerShiftReg_w1_d3_io_d),
    .io_q(SynchronizerShiftReg_w1_d3_io_q),
    .io_covSum(SynchronizerShiftReg_w1_d3_io_covSum),
    .metaAssert(SynchronizerShiftReg_w1_d3_metaAssert),
    .metaReset(SynchronizerShiftReg_w1_d3_metaReset)
  );
  assign auto_out_0 = SynchronizerShiftReg_w1_d3_io_q; // @[LazyModule.scala 173:49]
  assign SynchronizerShiftReg_w1_d3_clock = clock;
  assign SynchronizerShiftReg_w1_d3_io_d = auto_in_sync_0; // @[ShiftReg.scala 49:16]
  assign IntSyncCrossingSink_covSum = 30'h0;
  assign SynchronizerShiftReg_w1_d3_sum = IntSyncCrossingSink_covSum + SynchronizerShiftReg_w1_d3_io_covSum;
  assign io_covSum = SynchronizerShiftReg_w1_d3_sum;
  assign SynchronizerShiftReg_w1_d3_metaAssert_wire = SynchronizerShiftReg_w1_d3_metaAssert;
  assign metaAssert = SynchronizerShiftReg_w1_d3_metaAssert_wire;
  assign SynchronizerShiftReg_w1_d3_metaReset = metaReset | SynchronizerShiftReg_w1_d3_halt;
endmodule
module IntSyncCrossingSink_1(
  input         auto_in_sync_0,
  input         auto_in_sync_1,
  output        auto_out_0,
  output        auto_out_1,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [29:0] IntSyncCrossingSink_1_covSum;
  assign auto_out_0 = auto_in_sync_0; // @[LazyModule.scala 173:49]
  assign auto_out_1 = auto_in_sync_1; // @[LazyModule.scala 173:49]
  assign IntSyncCrossingSink_1_covSum = 30'h0;
  assign io_covSum = IntSyncCrossingSink_1_covSum;
  assign metaAssert = 1'h0;
endmodule
module IntSyncCrossingSink_2(
  input         auto_in_sync_0,
  output        auto_out_0,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [29:0] IntSyncCrossingSink_2_covSum;
  assign auto_out_0 = auto_in_sync_0; // @[LazyModule.scala 173:49]
  assign IntSyncCrossingSink_2_covSum = 30'h0;
  assign io_covSum = IntSyncCrossingSink_2_covSum;
  assign metaAssert = 1'h0;
endmodule
module FPU(
  input         clock,
  input         reset,
  input  [31:0] io_inst,
  input  [63:0] io_fromint_data,
  input  [2:0]  io_fcsr_rm,
  output        io_fcsr_flags_valid,
  output [4:0]  io_fcsr_flags_bits,
  output [63:0] io_store_data,
  output [63:0] io_toint_data,
  input         io_dmem_resp_val,
  input  [2:0]  io_dmem_resp_type,
  input  [4:0]  io_dmem_resp_tag,
  input  [63:0] io_dmem_resp_data,
  input         io_valid,
  output        io_fcsr_rdy,
  output        io_nack_mem,
  output        io_illegal_rm,
  input         io_killx,
  input         io_killm,
  output        io_dec_wen,
  output        io_dec_ren1,
  output        io_dec_ren2,
  output        io_dec_ren3,
  output        io_sboard_set,
  output        io_sboard_clr,
  output [4:0]  io_sboard_clra,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         dfma_halt,
  input         fpmu_halt,
  input         divSqrt_1_halt,
  input         ifpu_halt,
  input         divSqrt_halt,
  input         fpiu_halt,
  input         sfma_halt
);
  wire [31:0] fp_decoder_io_inst; // @[FPU.scala 674:26]
  wire  fp_decoder_io_sigs_wen; // @[FPU.scala 674:26]
  wire  fp_decoder_io_sigs_ren1; // @[FPU.scala 674:26]
  wire  fp_decoder_io_sigs_ren2; // @[FPU.scala 674:26]
  wire  fp_decoder_io_sigs_ren3; // @[FPU.scala 674:26]
  wire  fp_decoder_io_sigs_swap12; // @[FPU.scala 674:26]
  wire  fp_decoder_io_sigs_swap23; // @[FPU.scala 674:26]
  wire  fp_decoder_io_sigs_singleIn; // @[FPU.scala 674:26]
  wire  fp_decoder_io_sigs_singleOut; // @[FPU.scala 674:26]
  wire  fp_decoder_io_sigs_fromint; // @[FPU.scala 674:26]
  wire  fp_decoder_io_sigs_toint; // @[FPU.scala 674:26]
  wire  fp_decoder_io_sigs_fastpipe; // @[FPU.scala 674:26]
  wire  fp_decoder_io_sigs_fma; // @[FPU.scala 674:26]
  wire  fp_decoder_io_sigs_div; // @[FPU.scala 674:26]
  wire  fp_decoder_io_sigs_sqrt; // @[FPU.scala 674:26]
  wire  fp_decoder_io_sigs_wflags; // @[FPU.scala 674:26]
  wire [29:0] fp_decoder_io_covSum; // @[FPU.scala 674:26]
  wire  fp_decoder_metaAssert; // @[FPU.scala 674:26]
  reg [64:0] regfile [0:31]; // @[FPU.scala 715:20]
  reg [95:0] _RAND_0;
  wire [64:0] regfile__T_499_data; // @[FPU.scala 715:20]
  wire [4:0] regfile__T_499_addr; // @[FPU.scala 715:20]
  wire [64:0] regfile__T_502_data; // @[FPU.scala 715:20]
  wire [4:0] regfile__T_502_addr; // @[FPU.scala 715:20]
  wire [64:0] regfile__T_505_data; // @[FPU.scala 715:20]
  wire [4:0] regfile__T_505_addr; // @[FPU.scala 715:20]
  wire [64:0] regfile__T_472_data; // @[FPU.scala 715:20]
  wire [4:0] regfile__T_472_addr; // @[FPU.scala 715:20]
  wire  regfile__T_472_mask; // @[FPU.scala 715:20]
  wire  regfile__T_472_en; // @[FPU.scala 715:20]
  wire [64:0] regfile__T_1002_data; // @[FPU.scala 715:20]
  wire [4:0] regfile__T_1002_addr; // @[FPU.scala 715:20]
  wire  regfile__T_1002_mask; // @[FPU.scala 715:20]
  wire  regfile__T_1002_en; // @[FPU.scala 715:20]
  wire  sfma_clock; // @[FPU.scala 759:20]
  wire  sfma_reset; // @[FPU.scala 759:20]
  wire  sfma_io_in_valid; // @[FPU.scala 759:20]
  wire  sfma_io_in_bits_ren3; // @[FPU.scala 759:20]
  wire  sfma_io_in_bits_swap23; // @[FPU.scala 759:20]
  wire [2:0] sfma_io_in_bits_rm; // @[FPU.scala 759:20]
  wire [1:0] sfma_io_in_bits_fmaCmd; // @[FPU.scala 759:20]
  wire [64:0] sfma_io_in_bits_in1; // @[FPU.scala 759:20]
  wire [64:0] sfma_io_in_bits_in2; // @[FPU.scala 759:20]
  wire [64:0] sfma_io_in_bits_in3; // @[FPU.scala 759:20]
  wire [64:0] sfma_io_out_bits_data; // @[FPU.scala 759:20]
  wire [4:0] sfma_io_out_bits_exc; // @[FPU.scala 759:20]
  wire [29:0] sfma_io_covSum; // @[FPU.scala 759:20]
  wire  sfma_metaAssert; // @[FPU.scala 759:20]
  wire  sfma_metaReset; // @[FPU.scala 759:20]
  wire  sfma_fma_halt; // @[FPU.scala 759:20]
  wire  fpiu_clock; // @[FPU.scala 763:20]
  wire  fpiu_io_in_valid; // @[FPU.scala 763:20]
  wire  fpiu_io_in_bits_ren2; // @[FPU.scala 763:20]
  wire  fpiu_io_in_bits_singleIn; // @[FPU.scala 763:20]
  wire  fpiu_io_in_bits_singleOut; // @[FPU.scala 763:20]
  wire  fpiu_io_in_bits_wflags; // @[FPU.scala 763:20]
  wire [2:0] fpiu_io_in_bits_rm; // @[FPU.scala 763:20]
  wire [1:0] fpiu_io_in_bits_typ; // @[FPU.scala 763:20]
  wire [64:0] fpiu_io_in_bits_in1; // @[FPU.scala 763:20]
  wire [64:0] fpiu_io_in_bits_in2; // @[FPU.scala 763:20]
  wire [2:0] fpiu_io_out_bits_in_rm; // @[FPU.scala 763:20]
  wire [64:0] fpiu_io_out_bits_in_in1; // @[FPU.scala 763:20]
  wire [64:0] fpiu_io_out_bits_in_in2; // @[FPU.scala 763:20]
  wire  fpiu_io_out_bits_lt; // @[FPU.scala 763:20]
  wire [63:0] fpiu_io_out_bits_store; // @[FPU.scala 763:20]
  wire [63:0] fpiu_io_out_bits_toint; // @[FPU.scala 763:20]
  wire [4:0] fpiu_io_out_bits_exc; // @[FPU.scala 763:20]
  wire [29:0] fpiu_io_covSum; // @[FPU.scala 763:20]
  wire  fpiu_metaAssert; // @[FPU.scala 763:20]
  wire  fpiu_metaReset; // @[FPU.scala 763:20]
  wire  ifpu_clock; // @[FPU.scala 773:20]
  wire  ifpu_reset; // @[FPU.scala 773:20]
  wire  ifpu_io_in_valid; // @[FPU.scala 773:20]
  wire  ifpu_io_in_bits_singleIn; // @[FPU.scala 773:20]
  wire  ifpu_io_in_bits_wflags; // @[FPU.scala 773:20]
  wire [2:0] ifpu_io_in_bits_rm; // @[FPU.scala 773:20]
  wire [1:0] ifpu_io_in_bits_typ; // @[FPU.scala 773:20]
  wire [63:0] ifpu_io_in_bits_in1; // @[FPU.scala 773:20]
  wire [64:0] ifpu_io_out_bits_data; // @[FPU.scala 773:20]
  wire [4:0] ifpu_io_out_bits_exc; // @[FPU.scala 773:20]
  wire [29:0] ifpu_io_covSum; // @[FPU.scala 773:20]
  wire  ifpu_metaAssert; // @[FPU.scala 773:20]
  wire  ifpu_metaReset; // @[FPU.scala 773:20]
  wire  fpmu_clock; // @[FPU.scala 778:20]
  wire  fpmu_reset; // @[FPU.scala 778:20]
  wire  fpmu_io_in_valid; // @[FPU.scala 778:20]
  wire  fpmu_io_in_bits_ren2; // @[FPU.scala 778:20]
  wire  fpmu_io_in_bits_singleOut; // @[FPU.scala 778:20]
  wire  fpmu_io_in_bits_wflags; // @[FPU.scala 778:20]
  wire [2:0] fpmu_io_in_bits_rm; // @[FPU.scala 778:20]
  wire [64:0] fpmu_io_in_bits_in1; // @[FPU.scala 778:20]
  wire [64:0] fpmu_io_in_bits_in2; // @[FPU.scala 778:20]
  wire [64:0] fpmu_io_out_bits_data; // @[FPU.scala 778:20]
  wire [4:0] fpmu_io_out_bits_exc; // @[FPU.scala 778:20]
  wire  fpmu_io_lt; // @[FPU.scala 778:20]
  wire [29:0] fpmu_io_covSum; // @[FPU.scala 778:20]
  wire  fpmu_metaAssert; // @[FPU.scala 778:20]
  wire  fpmu_metaReset; // @[FPU.scala 778:20]
  wire  dfma_clock; // @[FPU.scala 797:28]
  wire  dfma_reset; // @[FPU.scala 797:28]
  wire  dfma_io_in_valid; // @[FPU.scala 797:28]
  wire  dfma_io_in_bits_ren3; // @[FPU.scala 797:28]
  wire  dfma_io_in_bits_swap23; // @[FPU.scala 797:28]
  wire [2:0] dfma_io_in_bits_rm; // @[FPU.scala 797:28]
  wire [1:0] dfma_io_in_bits_fmaCmd; // @[FPU.scala 797:28]
  wire [64:0] dfma_io_in_bits_in1; // @[FPU.scala 797:28]
  wire [64:0] dfma_io_in_bits_in2; // @[FPU.scala 797:28]
  wire [64:0] dfma_io_in_bits_in3; // @[FPU.scala 797:28]
  wire [64:0] dfma_io_out_bits_data; // @[FPU.scala 797:28]
  wire [4:0] dfma_io_out_bits_exc; // @[FPU.scala 797:28]
  wire [29:0] dfma_io_covSum; // @[FPU.scala 797:28]
  wire  dfma_metaAssert; // @[FPU.scala 797:28]
  wire  dfma_metaReset; // @[FPU.scala 797:28]
  wire  dfma_fma_halt; // @[FPU.scala 797:28]
  wire  divSqrt_clock; // @[FPU.scala 887:27]
  wire  divSqrt_reset; // @[FPU.scala 887:27]
  wire  divSqrt_io_inReady; // @[FPU.scala 887:27]
  wire  divSqrt_io_inValid; // @[FPU.scala 887:27]
  wire  divSqrt_io_sqrtOp; // @[FPU.scala 887:27]
  wire [32:0] divSqrt_io_a; // @[FPU.scala 887:27]
  wire [32:0] divSqrt_io_b; // @[FPU.scala 887:27]
  wire [2:0] divSqrt_io_roundingMode; // @[FPU.scala 887:27]
  wire  divSqrt_io_outValid_div; // @[FPU.scala 887:27]
  wire  divSqrt_io_outValid_sqrt; // @[FPU.scala 887:27]
  wire [32:0] divSqrt_io_out; // @[FPU.scala 887:27]
  wire [4:0] divSqrt_io_exceptionFlags; // @[FPU.scala 887:27]
  wire [29:0] divSqrt_io_covSum; // @[FPU.scala 887:27]
  wire  divSqrt_metaAssert; // @[FPU.scala 887:27]
  wire  divSqrt_metaReset; // @[FPU.scala 887:27]
  wire  divSqrt_divSqrtRecFNToRaw_halt; // @[FPU.scala 887:27]
  wire  divSqrt_1_clock; // @[FPU.scala 887:27]
  wire  divSqrt_1_reset; // @[FPU.scala 887:27]
  wire  divSqrt_1_io_inReady; // @[FPU.scala 887:27]
  wire  divSqrt_1_io_inValid; // @[FPU.scala 887:27]
  wire  divSqrt_1_io_sqrtOp; // @[FPU.scala 887:27]
  wire [64:0] divSqrt_1_io_a; // @[FPU.scala 887:27]
  wire [64:0] divSqrt_1_io_b; // @[FPU.scala 887:27]
  wire [2:0] divSqrt_1_io_roundingMode; // @[FPU.scala 887:27]
  wire  divSqrt_1_io_outValid_div; // @[FPU.scala 887:27]
  wire  divSqrt_1_io_outValid_sqrt; // @[FPU.scala 887:27]
  wire [64:0] divSqrt_1_io_out; // @[FPU.scala 887:27]
  wire [4:0] divSqrt_1_io_exceptionFlags; // @[FPU.scala 887:27]
  wire [29:0] divSqrt_1_io_covSum; // @[FPU.scala 887:27]
  wire  divSqrt_1_metaAssert; // @[FPU.scala 887:27]
  wire  divSqrt_1_metaReset; // @[FPU.scala 887:27]
  wire  divSqrt_1_divSqrtRecFNToRaw_halt; // @[FPU.scala 887:27]
  reg  ex_reg_valid; // @[FPU.scala 678:25]
  reg [31:0] _RAND_1;
  reg [31:0] ex_reg_inst; // @[Reg.scala 11:16]
  reg [31:0] _RAND_2;
  reg  ex_reg_ctrl_ren2; // @[Reg.scala 11:16]
  reg [31:0] _RAND_3;
  reg  ex_reg_ctrl_ren3; // @[Reg.scala 11:16]
  reg [31:0] _RAND_4;
  reg  ex_reg_ctrl_swap23; // @[Reg.scala 11:16]
  reg [31:0] _RAND_5;
  reg  ex_reg_ctrl_singleIn; // @[Reg.scala 11:16]
  reg [31:0] _RAND_6;
  reg  ex_reg_ctrl_singleOut; // @[Reg.scala 11:16]
  reg [31:0] _RAND_7;
  reg  ex_reg_ctrl_fromint; // @[Reg.scala 11:16]
  reg [31:0] _RAND_8;
  reg  ex_reg_ctrl_toint; // @[Reg.scala 11:16]
  reg [31:0] _RAND_9;
  reg  ex_reg_ctrl_fastpipe; // @[Reg.scala 11:16]
  reg [31:0] _RAND_10;
  reg  ex_reg_ctrl_fma; // @[Reg.scala 11:16]
  reg [31:0] _RAND_11;
  reg  ex_reg_ctrl_div; // @[Reg.scala 11:16]
  reg [31:0] _RAND_12;
  reg  ex_reg_ctrl_sqrt; // @[Reg.scala 11:16]
  reg [31:0] _RAND_13;
  reg  ex_reg_ctrl_wflags; // @[Reg.scala 11:16]
  reg [31:0] _RAND_14;
  reg [4:0] ex_ra_0; // @[FPU.scala 681:31]
  reg [31:0] _RAND_15;
  reg [4:0] ex_ra_1; // @[FPU.scala 681:31]
  reg [31:0] _RAND_16;
  reg [4:0] ex_ra_2; // @[FPU.scala 681:31]
  reg [31:0] _RAND_17;
  reg  mem_reg_valid; // @[FPU.scala 689:30]
  reg [31:0] _RAND_18;
  wire  killm; // @[FPU.scala 690:25]
  wire  _T_47; // @[FPU.scala 694:41]
  wire  killx; // @[FPU.scala 694:24]
  wire  _T_49; // @[FPU.scala 695:33]
  reg [31:0] mem_reg_inst; // @[Reg.scala 11:16]
  reg [31:0] _RAND_19;
  wire  _T_54; // @[FPU.scala 697:45]
  reg  wb_reg_valid; // @[FPU.scala 697:25]
  reg [31:0] _RAND_20;
  reg  mem_ctrl_singleOut; // @[Reg.scala 11:16]
  reg [31:0] _RAND_21;
  reg  mem_ctrl_fromint; // @[Reg.scala 11:16]
  reg [31:0] _RAND_22;
  reg  mem_ctrl_toint; // @[Reg.scala 11:16]
  reg [31:0] _RAND_23;
  reg  mem_ctrl_fastpipe; // @[Reg.scala 11:16]
  reg [31:0] _RAND_24;
  reg  mem_ctrl_fma; // @[Reg.scala 11:16]
  reg [31:0] _RAND_25;
  reg  mem_ctrl_div; // @[Reg.scala 11:16]
  reg [31:0] _RAND_26;
  reg  mem_ctrl_sqrt; // @[Reg.scala 11:16]
  reg [31:0] _RAND_27;
  reg  mem_ctrl_wflags; // @[Reg.scala 11:16]
  reg [31:0] _RAND_28;
  reg  wb_ctrl_toint; // @[Reg.scala 11:16]
  reg [31:0] _RAND_29;
  reg  load_wb; // @[FPU.scala 709:20]
  reg [31:0] _RAND_30;
  reg  load_wb_double; // @[Reg.scala 11:16]
  reg [31:0] _RAND_31;
  reg [63:0] load_wb_data; // @[Reg.scala 11:16]
  reg [63:0] _RAND_32;
  reg [4:0] load_wb_tag; // @[Reg.scala 11:16]
  reg [31:0] _RAND_33;
  wire [63:0] _T_67; // @[package.scala 31:71]
  wire [63:0] _T_68; // @[FPU.scala 358:23]
  wire  _T_72; // @[rawFloatFromFN.scala 50:34]
  wire  _T_73; // @[rawFloatFromFN.scala 51:38]
  wire [31:0] _T_78; // @[Bitwise.scala 103:31]
  wire [31:0] _T_80; // @[Bitwise.scala 103:65]
  wire [31:0] _T_82; // @[Bitwise.scala 103:75]
  wire [31:0] _T_83; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_165; // @[Bitwise.scala 103:31]
  wire [31:0] _T_88; // @[Bitwise.scala 103:31]
  wire [31:0] _T_90; // @[Bitwise.scala 103:65]
  wire [31:0] _T_92; // @[Bitwise.scala 103:75]
  wire [31:0] _T_93; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_166; // @[Bitwise.scala 103:31]
  wire [31:0] _T_98; // @[Bitwise.scala 103:31]
  wire [31:0] _T_100; // @[Bitwise.scala 103:65]
  wire [31:0] _T_102; // @[Bitwise.scala 103:75]
  wire [31:0] _T_103; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_167; // @[Bitwise.scala 103:31]
  wire [31:0] _T_108; // @[Bitwise.scala 103:31]
  wire [31:0] _T_110; // @[Bitwise.scala 103:65]
  wire [31:0] _T_112; // @[Bitwise.scala 103:75]
  wire [31:0] _T_113; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_168; // @[Bitwise.scala 103:31]
  wire [31:0] _T_118; // @[Bitwise.scala 103:31]
  wire [31:0] _T_120; // @[Bitwise.scala 103:65]
  wire [31:0] _T_122; // @[Bitwise.scala 103:75]
  wire [31:0] _T_123; // @[Bitwise.scala 103:39]
  wire [15:0] _T_129; // @[Bitwise.scala 103:31]
  wire [15:0] _T_131; // @[Bitwise.scala 103:65]
  wire [15:0] _T_133; // @[Bitwise.scala 103:75]
  wire [15:0] _T_134; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_169; // @[Bitwise.scala 103:31]
  wire [15:0] _T_139; // @[Bitwise.scala 103:31]
  wire [15:0] _T_141; // @[Bitwise.scala 103:65]
  wire [15:0] _T_143; // @[Bitwise.scala 103:75]
  wire [15:0] _T_144; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_170; // @[Bitwise.scala 103:31]
  wire [15:0] _T_149; // @[Bitwise.scala 103:31]
  wire [15:0] _T_151; // @[Bitwise.scala 103:65]
  wire [15:0] _T_153; // @[Bitwise.scala 103:75]
  wire [15:0] _T_154; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_171; // @[Bitwise.scala 103:31]
  wire [15:0] _T_159; // @[Bitwise.scala 103:31]
  wire [15:0] _T_161; // @[Bitwise.scala 103:65]
  wire [15:0] _T_163; // @[Bitwise.scala 103:75]
  wire [15:0] _T_164; // @[Bitwise.scala 103:39]
  wire [51:0] _T_176; // @[Cat.scala 30:58]
  wire [5:0] _T_229; // @[Mux.scala 31:69]
  wire [5:0] _T_230; // @[Mux.scala 31:69]
  wire [5:0] _T_231; // @[Mux.scala 31:69]
  wire [5:0] _T_232; // @[Mux.scala 31:69]
  wire [5:0] _T_233; // @[Mux.scala 31:69]
  wire [5:0] _T_234; // @[Mux.scala 31:69]
  wire [5:0] _T_235; // @[Mux.scala 31:69]
  wire [5:0] _T_236; // @[Mux.scala 31:69]
  wire [5:0] _T_237; // @[Mux.scala 31:69]
  wire [5:0] _T_238; // @[Mux.scala 31:69]
  wire [5:0] _T_239; // @[Mux.scala 31:69]
  wire [5:0] _T_240; // @[Mux.scala 31:69]
  wire [5:0] _T_241; // @[Mux.scala 31:69]
  wire [5:0] _T_242; // @[Mux.scala 31:69]
  wire [5:0] _T_243; // @[Mux.scala 31:69]
  wire [5:0] _T_244; // @[Mux.scala 31:69]
  wire [5:0] _T_245; // @[Mux.scala 31:69]
  wire [5:0] _T_246; // @[Mux.scala 31:69]
  wire [5:0] _T_247; // @[Mux.scala 31:69]
  wire [5:0] _T_248; // @[Mux.scala 31:69]
  wire [5:0] _T_249; // @[Mux.scala 31:69]
  wire [5:0] _T_250; // @[Mux.scala 31:69]
  wire [5:0] _T_251; // @[Mux.scala 31:69]
  wire [5:0] _T_252; // @[Mux.scala 31:69]
  wire [5:0] _T_253; // @[Mux.scala 31:69]
  wire [5:0] _T_254; // @[Mux.scala 31:69]
  wire [5:0] _T_255; // @[Mux.scala 31:69]
  wire [5:0] _T_256; // @[Mux.scala 31:69]
  wire [5:0] _T_257; // @[Mux.scala 31:69]
  wire [5:0] _T_258; // @[Mux.scala 31:69]
  wire [5:0] _T_259; // @[Mux.scala 31:69]
  wire [5:0] _T_260; // @[Mux.scala 31:69]
  wire [5:0] _T_261; // @[Mux.scala 31:69]
  wire [5:0] _T_262; // @[Mux.scala 31:69]
  wire [5:0] _T_263; // @[Mux.scala 31:69]
  wire [5:0] _T_264; // @[Mux.scala 31:69]
  wire [5:0] _T_265; // @[Mux.scala 31:69]
  wire [5:0] _T_266; // @[Mux.scala 31:69]
  wire [5:0] _T_267; // @[Mux.scala 31:69]
  wire [5:0] _T_268; // @[Mux.scala 31:69]
  wire [5:0] _T_269; // @[Mux.scala 31:69]
  wire [5:0] _T_270; // @[Mux.scala 31:69]
  wire [5:0] _T_271; // @[Mux.scala 31:69]
  wire [5:0] _T_272; // @[Mux.scala 31:69]
  wire [5:0] _T_273; // @[Mux.scala 31:69]
  wire [5:0] _T_274; // @[Mux.scala 31:69]
  wire [5:0] _T_275; // @[Mux.scala 31:69]
  wire [5:0] _T_276; // @[Mux.scala 31:69]
  wire [5:0] _T_277; // @[Mux.scala 31:69]
  wire [5:0] _T_278; // @[Mux.scala 31:69]
  wire [5:0] _T_279; // @[Mux.scala 31:69]
  wire [114:0] _GEN_172; // @[rawFloatFromFN.scala 54:36]
  wire [114:0] _T_280; // @[rawFloatFromFN.scala 54:36]
  wire [51:0] _T_282; // @[rawFloatFromFN.scala 54:64]
  wire [11:0] _GEN_173; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_283; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_284; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_285; // @[rawFloatFromFN.scala 60:27]
  wire [10:0] _GEN_174; // @[rawFloatFromFN.scala 60:22]
  wire [10:0] _T_286; // @[rawFloatFromFN.scala 60:22]
  wire [11:0] _GEN_175; // @[rawFloatFromFN.scala 59:15]
  wire [11:0] _T_288; // @[rawFloatFromFN.scala 59:15]
  wire  _T_289; // @[rawFloatFromFN.scala 62:34]
  wire  _T_291; // @[rawFloatFromFN.scala 63:62]
  wire  _T_295; // @[rawFloatFromFN.scala 66:33]
  wire [12:0] _T_298; // @[rawFloatFromFN.scala 70:48]
  wire [51:0] _T_300; // @[rawFloatFromFN.scala 72:42]
  wire [53:0] _T_302; // @[Cat.scala 30:58]
  wire [2:0] _T_304; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_176; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_306; // @[recFNFromFN.scala 48:79]
  wire [64:0] _T_311; // @[Cat.scala 30:58]
  wire  _T_315; // @[rawFloatFromFN.scala 50:34]
  wire  _T_316; // @[rawFloatFromFN.scala 51:38]
  wire [15:0] _T_321; // @[Bitwise.scala 103:31]
  wire [15:0] _T_323; // @[Bitwise.scala 103:65]
  wire [15:0] _T_325; // @[Bitwise.scala 103:75]
  wire [15:0] _T_326; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_177; // @[Bitwise.scala 103:31]
  wire [15:0] _T_331; // @[Bitwise.scala 103:31]
  wire [15:0] _T_333; // @[Bitwise.scala 103:65]
  wire [15:0] _T_335; // @[Bitwise.scala 103:75]
  wire [15:0] _T_336; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_178; // @[Bitwise.scala 103:31]
  wire [15:0] _T_341; // @[Bitwise.scala 103:31]
  wire [15:0] _T_343; // @[Bitwise.scala 103:65]
  wire [15:0] _T_345; // @[Bitwise.scala 103:75]
  wire [15:0] _T_346; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_179; // @[Bitwise.scala 103:31]
  wire [15:0] _T_351; // @[Bitwise.scala 103:31]
  wire [15:0] _T_353; // @[Bitwise.scala 103:65]
  wire [15:0] _T_355; // @[Bitwise.scala 103:75]
  wire [15:0] _T_356; // @[Bitwise.scala 103:39]
  wire [22:0] _T_376; // @[Cat.scala 30:58]
  wire [4:0] _T_400; // @[Mux.scala 31:69]
  wire [4:0] _T_401; // @[Mux.scala 31:69]
  wire [4:0] _T_402; // @[Mux.scala 31:69]
  wire [4:0] _T_403; // @[Mux.scala 31:69]
  wire [4:0] _T_404; // @[Mux.scala 31:69]
  wire [4:0] _T_405; // @[Mux.scala 31:69]
  wire [4:0] _T_406; // @[Mux.scala 31:69]
  wire [4:0] _T_407; // @[Mux.scala 31:69]
  wire [4:0] _T_408; // @[Mux.scala 31:69]
  wire [4:0] _T_409; // @[Mux.scala 31:69]
  wire [4:0] _T_410; // @[Mux.scala 31:69]
  wire [4:0] _T_411; // @[Mux.scala 31:69]
  wire [4:0] _T_412; // @[Mux.scala 31:69]
  wire [4:0] _T_413; // @[Mux.scala 31:69]
  wire [4:0] _T_414; // @[Mux.scala 31:69]
  wire [4:0] _T_415; // @[Mux.scala 31:69]
  wire [4:0] _T_416; // @[Mux.scala 31:69]
  wire [4:0] _T_417; // @[Mux.scala 31:69]
  wire [4:0] _T_418; // @[Mux.scala 31:69]
  wire [4:0] _T_419; // @[Mux.scala 31:69]
  wire [4:0] _T_420; // @[Mux.scala 31:69]
  wire [4:0] _T_421; // @[Mux.scala 31:69]
  wire [53:0] _GEN_180; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_422; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_424; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_181; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_425; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_426; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_427; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_182; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_428; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_183; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_430; // @[rawFloatFromFN.scala 59:15]
  wire  _T_431; // @[rawFloatFromFN.scala 62:34]
  wire  _T_433; // @[rawFloatFromFN.scala 63:62]
  wire  _T_437; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_440; // @[rawFloatFromFN.scala 70:48]
  wire [22:0] _T_442; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_444; // @[Cat.scala 30:58]
  wire [2:0] _T_446; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_184; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_448; // @[recFNFromFN.scala 48:79]
  wire [32:0] _T_453; // @[Cat.scala 30:58]
  wire  _T_457; // @[FPU.scala 265:42]
  wire [64:0] _T_468; // @[Cat.scala 30:58]
  wire  _T_471; // @[FPU.scala 197:56]
  wire [64:0] wdata; // @[FPU.scala 271:8]
  wire  _T_485; // @[FPU.scala 197:56]
  wire  _T_490; // @[FPU.scala 312:96]
  wire  _T_491; // @[FPU.scala 312:55]
  wire  _T_492; // @[FPU.scala 312:31]
  wire  _T_495; // @[FPU.scala 719:11]
  wire  _T_513; // @[FPU.scala 733:29]
  wire  _T_517; // @[FPU.scala 737:38]
  wire  _T_519; // @[FPU.scala 760:33]
  wire  tag; // @[FPU.scala 741:15]
  wire [32:0] _T_526; // @[Cat.scala 30:58]
  wire  _T_529; // @[FPU.scala 259:84]
  wire [32:0] _T_551; // @[FPU.scala 299:31]
  wire [32:0] _T_552; // @[FPU.scala 299:26]
  wire [32:0] _T_557; // @[Cat.scala 30:58]
  wire  _T_560; // @[FPU.scala 259:84]
  wire [32:0] _T_582; // @[FPU.scala 299:31]
  wire [32:0] _T_583; // @[FPU.scala 299:26]
  wire [32:0] _T_588; // @[Cat.scala 30:58]
  wire  _T_591; // @[FPU.scala 259:84]
  wire [32:0] _T_613; // @[FPU.scala 299:31]
  wire [32:0] _T_614; // @[FPU.scala 299:26]
  wire  _T_619; // @[FPU.scala 748:53]
  wire [1:0] _GEN_185; // @[FPU.scala 748:36]
  wire  _T_621; // @[FPU.scala 764:51]
  wire  _T_622; // @[FPU.scala 764:66]
  wire  _T_623; // @[FPU.scala 764:103]
  wire  _T_624; // @[FPU.scala 764:82]
  wire [75:0] _T_635; // @[FPU.scala 225:28]
  wire [11:0] _GEN_186; // @[FPU.scala 228:31]
  wire [11:0] _T_639; // @[FPU.scala 228:31]
  wire [11:0] _T_642; // @[FPU.scala 228:48]
  wire  _T_643; // @[FPU.scala 229:19]
  wire  _T_644; // @[FPU.scala 229:36]
  wire  _T_645; // @[FPU.scala 229:25]
  wire [11:0] _T_647; // @[Cat.scala 30:58]
  wire [11:0] _T_649; // @[FPU.scala 229:10]
  wire [64:0] _T_651; // @[Cat.scala 30:58]
  wire  _T_657; // @[package.scala 31:71]
  wire [64:0] _T_659; // @[package.scala 31:71]
  wire [75:0] _T_669; // @[FPU.scala 225:28]
  wire [11:0] _GEN_187; // @[FPU.scala 228:31]
  wire [11:0] _T_673; // @[FPU.scala 228:31]
  wire [11:0] _T_676; // @[FPU.scala 228:48]
  wire  _T_677; // @[FPU.scala 229:19]
  wire  _T_678; // @[FPU.scala 229:36]
  wire  _T_679; // @[FPU.scala 229:25]
  wire [11:0] _T_681; // @[Cat.scala 30:58]
  wire [11:0] _T_683; // @[FPU.scala 229:10]
  wire [64:0] _T_685; // @[Cat.scala 30:58]
  wire  _T_691; // @[package.scala 31:71]
  wire [64:0] _T_693; // @[package.scala 31:71]
  wire [64:0] _T_738; // @[FPU.scala 776:29]
  reg [4:0] divSqrt_waddr; // @[FPU.scala 785:26]
  reg [31:0] _RAND_34;
  wire  _T_851; // @[FPU.scala 795:56]
  wire [1:0] _T_852; // @[FPU.scala 804:23]
  wire  _T_854; // @[FPU.scala 800:62]
  wire [2:0] _T_855; // @[FPU.scala 804:23]
  wire  _T_856; // @[FPU.scala 804:78]
  wire [1:0] _GEN_194; // @[FPU.scala 804:78]
  wire [1:0] _T_857; // @[FPU.scala 804:78]
  wire [2:0] _GEN_195; // @[FPU.scala 804:78]
  wire [2:0] memLatencyMask; // @[FPU.scala 804:78]
  reg [2:0] wen; // @[FPU.scala 818:16]
  reg [31:0] _RAND_35;
  reg [4:0] wbInfo_0_rd; // @[FPU.scala 819:19]
  reg [31:0] _RAND_36;
  reg  wbInfo_0_single; // @[FPU.scala 819:19]
  reg [31:0] _RAND_37;
  reg [1:0] wbInfo_0_pipeid; // @[FPU.scala 819:19]
  reg [31:0] _RAND_38;
  reg [4:0] wbInfo_1_rd; // @[FPU.scala 819:19]
  reg [31:0] _RAND_39;
  reg  wbInfo_1_single; // @[FPU.scala 819:19]
  reg [31:0] _RAND_40;
  reg [1:0] wbInfo_1_pipeid; // @[FPU.scala 819:19]
  reg [31:0] _RAND_41;
  reg [4:0] wbInfo_2_rd; // @[FPU.scala 819:19]
  reg [31:0] _RAND_42;
  reg  wbInfo_2_single; // @[FPU.scala 819:19]
  reg [31:0] _RAND_43;
  reg [1:0] wbInfo_2_pipeid; // @[FPU.scala 819:19]
  reg [31:0] _RAND_44;
  wire  _T_867; // @[FPU.scala 820:48]
  wire  _T_868; // @[FPU.scala 820:69]
  wire  mem_wen; // @[FPU.scala 820:31]
  wire [1:0] _T_869; // @[FPU.scala 804:23]
  wire [1:0] _T_870; // @[FPU.scala 804:23]
  wire  _T_871; // @[FPU.scala 795:56]
  wire [2:0] _T_872; // @[FPU.scala 804:23]
  wire  _T_874; // @[FPU.scala 800:62]
  wire [3:0] _T_875; // @[FPU.scala 804:23]
  wire [1:0] _T_876; // @[FPU.scala 804:78]
  wire [2:0] _GEN_196; // @[FPU.scala 804:78]
  wire [2:0] _T_877; // @[FPU.scala 804:78]
  wire [3:0] _GEN_197; // @[FPU.scala 804:78]
  wire [3:0] _T_878; // @[FPU.scala 804:78]
  wire [3:0] _GEN_198; // @[FPU.scala 821:62]
  wire [3:0] _T_879; // @[FPU.scala 821:62]
  wire  _T_880; // @[FPU.scala 821:89]
  wire  _T_881; // @[FPU.scala 821:43]
  wire [2:0] _T_882; // @[FPU.scala 804:23]
  wire [2:0] _T_883; // @[FPU.scala 804:23]
  wire [3:0] _T_885; // @[FPU.scala 804:23]
  wire [4:0] _T_888; // @[FPU.scala 804:23]
  wire [2:0] _T_889; // @[FPU.scala 804:78]
  wire [3:0] _GEN_199; // @[FPU.scala 804:78]
  wire [3:0] _T_890; // @[FPU.scala 804:78]
  wire [4:0] _GEN_200; // @[FPU.scala 804:78]
  wire [4:0] _T_891; // @[FPU.scala 804:78]
  wire [4:0] _GEN_201; // @[FPU.scala 821:101]
  wire [4:0] _T_892; // @[FPU.scala 821:101]
  wire  _T_893; // @[FPU.scala 821:128]
  wire  _T_894; // @[FPU.scala 821:93]
  reg  write_port_busy; // @[Reg.scala 11:16]
  reg [31:0] _RAND_45;
  wire [2:0] _GEN_202; // @[FPU.scala 830:23]
  wire [2:0] _T_902; // @[FPU.scala 830:23]
  wire  _T_905; // @[FPU.scala 833:30]
  wire [1:0] _T_912; // @[FPU.scala 806:63]
  wire [1:0] _GEN_203; // @[FPU.scala 806:108]
  wire [1:0] _T_914; // @[FPU.scala 806:108]
  wire [1:0] _T_915; // @[FPU.scala 806:108]
  wire  _T_919; // @[FPU.scala 833:30]
  wire  _T_933; // @[FPU.scala 833:30]
  wire  divSqrt_typeTag; // @[FPU.scala 902:37]
  reg  divSqrt_killed; // @[FPU.scala 880:29]
  reg [31:0] _RAND_46;
  wire  _T_1111; // @[FPU.scala 902:37]
  wire  _GEN_154; // @[FPU.scala 902:66]
  wire  divSqrt_wen; // @[FPU.scala 902:66]
  wire  wdouble; // @[FPU.scala 843:20]
  wire  _T_946; // @[package.scala 31:81]
  wire [64:0] _T_947; // @[package.scala 31:71]
  wire  _T_948; // @[package.scala 31:81]
  wire [64:0] _T_949; // @[package.scala 31:71]
  wire  _T_950; // @[package.scala 31:81]
  wire [64:0] _T_951; // @[package.scala 31:71]
  wire  _T_1128; // @[FPU.scala 197:56]
  wire [64:0] _T_1125; // @[FPU.scala 340:25]
  wire [64:0] _T_1129; // @[FPU.scala 341:10]
  wire [32:0] _GEN_155; // @[FPU.scala 902:66]
  wire [64:0] divSqrt_wdata; // @[FPU.scala 902:66]
  wire [64:0] _T_952; // @[FPU.scala 844:22]
  wire [64:0] _T_963; // @[Cat.scala 30:58]
  wire [64:0] wdata_1; // @[package.scala 31:71]
  wire [4:0] _T_970; // @[package.scala 31:71]
  wire [4:0] _T_972; // @[package.scala 31:71]
  wire [4:0] wexc; // @[package.scala 31:71]
  wire  _T_977; // @[FPU.scala 846:35]
  wire  _T_990; // @[FPU.scala 197:56]
  wire  _T_995; // @[FPU.scala 312:96]
  wire  _T_996; // @[FPU.scala 312:55]
  wire  _T_997; // @[FPU.scala 312:31]
  wire  _T_1000; // @[FPU.scala 847:11]
  wire  wb_toint_valid; // @[FPU.scala 859:37]
  reg [4:0] wb_toint_exc; // @[Reg.scala 11:16]
  reg [31:0] _RAND_47;
  wire  _T_1007; // @[FPU.scala 861:41]
  wire [4:0] _T_1010; // @[FPU.scala 863:8]
  wire [4:0] _GEN_156; // @[FPU.scala 902:66]
  wire [4:0] divSqrt_flags; // @[FPU.scala 902:66]
  wire [4:0] _T_1011; // @[FPU.scala 864:8]
  wire [4:0] _T_1012; // @[FPU.scala 863:48]
  wire [4:0] _T_1014; // @[FPU.scala 865:8]
  wire  _T_1016; // @[FPU.scala 867:47]
  wire  _T_1017; // @[FPU.scala 867:72]
  wire  divSqrt_write_port_busy; // @[FPU.scala 867:65]
  wire  _T_1018; // @[FPU.scala 868:33]
  wire  _T_1019; // @[FPU.scala 868:68]
  wire  _T_1020; // @[FPU.scala 868:51]
  wire  _T_1022; // @[FPU.scala 868:87]
  wire  _T_1024; // @[FPU.scala 868:120]
  wire  divSqrt_inFlight; // @[FPU.scala 895:34]
  wire  _T_1025; // @[FPU.scala 868:131]
  wire  _T_1027; // @[FPU.scala 869:34]
  wire  _T_1034; // @[FPU.scala 872:96]
  reg  _T_1037; // @[FPU.scala 872:55]
  reg [31:0] _RAND_48;
  wire  _T_1043; // @[FPU.scala 873:60]
  wire  _T_1048; // @[package.scala 14:47]
  wire  _T_1049; // @[package.scala 14:47]
  wire  _T_1050; // @[package.scala 14:62]
  wire  _T_1052; // @[FPU.scala 877:67]
  wire  _T_1053; // @[FPU.scala 877:87]
  wire  _T_1054; // @[FPU.scala 877:73]
  wire  _T_1063; // @[FPU.scala 888:43]
  wire  _T_1065; // @[FPU.scala 888:65]
  wire [75:0] _T_1071; // @[FPU.scala 225:28]
  wire [11:0] _T_1075; // @[FPU.scala 228:31]
  wire [11:0] _T_1078; // @[FPU.scala 228:48]
  wire  _T_1079; // @[FPU.scala 229:19]
  wire  _T_1080; // @[FPU.scala 229:36]
  wire  _T_1081; // @[FPU.scala 229:25]
  wire [8:0] _T_1083; // @[Cat.scala 30:58]
  wire [8:0] _T_1085; // @[FPU.scala 229:10]
  wire [9:0] _T_1086; // @[Cat.scala 30:58]
  wire [75:0] _T_1091; // @[FPU.scala 225:28]
  wire [11:0] _T_1095; // @[FPU.scala 228:31]
  wire [11:0] _T_1098; // @[FPU.scala 228:48]
  wire  _T_1099; // @[FPU.scala 229:19]
  wire  _T_1100; // @[FPU.scala 229:36]
  wire  _T_1101; // @[FPU.scala 229:25]
  wire [8:0] _T_1103; // @[Cat.scala 30:58]
  wire [8:0] _T_1105; // @[FPU.scala 229:10]
  wire [9:0] _T_1106; // @[Cat.scala 30:58]
  wire  _T_1109; // @[FPU.scala 897:32]
  wire  _T_1114; // @[FPU.scala 888:43]
  wire  _T_1116; // @[FPU.scala 888:65]
  wire  _T_1120; // @[FPU.scala 897:32]
  reg [19:0] FPU_state; // @[Register tracking FPU state]
  reg [31:0] _RAND_49;
  reg  FPU_cov [0:1048575]; // @[Coverage map for FPU]
  reg [31:0] _RAND_50;
  wire  FPU_cov_read_data; // @[Coverage map for FPU]
  wire [19:0] FPU_cov_read_addr; // @[Coverage map for FPU]
  wire  FPU_cov_write_data; // @[Coverage map for FPU]
  wire [19:0] FPU_cov_write_addr; // @[Coverage map for FPU]
  wire  FPU_cov_write_mask; // @[Coverage map for FPU]
  wire  FPU_cov_write_en; // @[Coverage map for FPU]
  reg [29:0] FPU_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_51;
  wire [16:0] wen_shl;
  wire [19:0] wen_pad;
  wire [16:0] wb_reg_valid_shl;
  wire [19:0] wb_reg_valid_pad;
  wire [18:0] ex_reg_valid_shl;
  wire [19:0] ex_reg_valid_pad;
  wire [7:0] mem_ctrl_fma_shl;
  wire [19:0] mem_ctrl_fma_pad;
  wire [14:0] mem_ctrl_fromint_shl;
  wire [19:0] mem_ctrl_fromint_pad;
  wire [16:0] wbInfo_0_pipeid_shl;
  wire [19:0] wbInfo_0_pipeid_pad;
  wire [3:0] ex_reg_ctrl_fma_shl;
  wire [19:0] ex_reg_ctrl_fma_pad;
  wire [19:0] mem_reg_valid_shl;
  wire [19:0] mem_reg_valid_pad;
  wire [15:0] ex_reg_ctrl_singleIn_shl;
  wire [19:0] ex_reg_ctrl_singleIn_pad;
  wire [1:0] wbInfo_0_single_shl;
  wire [19:0] wbInfo_0_single_pad;
  wire [14:0] mem_ctrl_singleOut_shl;
  wire [19:0] mem_ctrl_singleOut_pad;
  wire [11:0] ex_reg_ctrl_singleOut_shl;
  wire [19:0] ex_reg_ctrl_singleOut_pad;
  wire [18:0] mem_ctrl_toint_shl;
  wire [19:0] mem_ctrl_toint_pad;
  wire [6:0] ex_reg_ctrl_fromint_shl;
  wire [19:0] ex_reg_ctrl_fromint_pad;
  wire [8:0] ex_reg_ctrl_fastpipe_shl;
  wire [19:0] ex_reg_ctrl_fastpipe_pad;
  wire [6:0] mem_ctrl_fastpipe_shl;
  wire [19:0] mem_ctrl_fastpipe_pad;
  wire [9:0] write_port_busy_shl;
  wire [19:0] write_port_busy_pad;
  wire [4:0] load_wb_double_shl;
  wire [19:0] load_wb_double_pad;
  wire [10:0] divSqrt_killed_shl;
  wire [19:0] divSqrt_killed_pad;
  wire [2:0] wb_ctrl_toint_shl;
  wire [19:0] wb_ctrl_toint_pad;
  wire [19:0] FPU_xor7;
  wire [19:0] FPU_xor18;
  wire [19:0] FPU_xor8;
  wire [19:0] FPU_xor3;
  wire [19:0] FPU_xor9;
  wire [19:0] FPU_xor22;
  wire [19:0] FPU_xor10;
  wire [19:0] FPU_xor4;
  wire [19:0] FPU_xor1;
  wire [19:0] FPU_xor11;
  wire [19:0] FPU_xor26;
  wire [19:0] FPU_xor12;
  wire [19:0] FPU_xor5;
  wire [19:0] FPU_xor13;
  wire [19:0] FPU_xor30;
  wire [19:0] FPU_xor14;
  wire [19:0] FPU_xor6;
  wire [19:0] FPU_xor2;
  wire [19:0] FPU_xor0;
  wire [29:0] fp_decoder_sum;
  wire [29:0] dfma_sum;
  wire [29:0] fpmu_sum;
  wire [29:0] divSqrt_1_sum;
  wire [29:0] ifpu_sum;
  wire [29:0] divSqrt_sum;
  wire [29:0] fpiu_sum;
  wire [29:0] sfma_sum;
  wire  stopEn0;
  wire  stopEn1;
  wire  ifpu_metaAssert_wire;
  wire  fpmu_metaAssert_wire;
  wire  fp_decoder_metaAssert_wire;
  wire  fpiu_metaAssert_wire;
  wire  divSqrt_1_metaAssert_wire;
  wire  divSqrt_metaAssert_wire;
  wire  dfma_metaAssert_wire;
  wire  sfma_metaAssert_wire;
  wire  FPU_or3;
  wire  FPU_or10;
  wire  FPU_or4;
  wire  FPU_or1;
  wire  FPU_or5;
  wire  FPU_or14;
  wire  FPU_or6;
  wire  FPU_or2;
  wire  FPU_or0;
  reg  FPU_metaAssert;
  reg [31:0] _RAND_52;
  FPUDecoder fp_decoder ( // @[FPU.scala 674:26]
    .io_inst(fp_decoder_io_inst),
    .io_sigs_wen(fp_decoder_io_sigs_wen),
    .io_sigs_ren1(fp_decoder_io_sigs_ren1),
    .io_sigs_ren2(fp_decoder_io_sigs_ren2),
    .io_sigs_ren3(fp_decoder_io_sigs_ren3),
    .io_sigs_swap12(fp_decoder_io_sigs_swap12),
    .io_sigs_swap23(fp_decoder_io_sigs_swap23),
    .io_sigs_singleIn(fp_decoder_io_sigs_singleIn),
    .io_sigs_singleOut(fp_decoder_io_sigs_singleOut),
    .io_sigs_fromint(fp_decoder_io_sigs_fromint),
    .io_sigs_toint(fp_decoder_io_sigs_toint),
    .io_sigs_fastpipe(fp_decoder_io_sigs_fastpipe),
    .io_sigs_fma(fp_decoder_io_sigs_fma),
    .io_sigs_div(fp_decoder_io_sigs_div),
    .io_sigs_sqrt(fp_decoder_io_sigs_sqrt),
    .io_sigs_wflags(fp_decoder_io_sigs_wflags),
    .io_covSum(fp_decoder_io_covSum),
    .metaAssert(fp_decoder_metaAssert)
  );
  FPUFMAPipe sfma ( // @[FPU.scala 759:20]
    .clock(sfma_clock),
    .reset(sfma_reset),
    .io_in_valid(sfma_io_in_valid),
    .io_in_bits_ren3(sfma_io_in_bits_ren3),
    .io_in_bits_swap23(sfma_io_in_bits_swap23),
    .io_in_bits_rm(sfma_io_in_bits_rm),
    .io_in_bits_fmaCmd(sfma_io_in_bits_fmaCmd),
    .io_in_bits_in1(sfma_io_in_bits_in1),
    .io_in_bits_in2(sfma_io_in_bits_in2),
    .io_in_bits_in3(sfma_io_in_bits_in3),
    .io_out_bits_data(sfma_io_out_bits_data),
    .io_out_bits_exc(sfma_io_out_bits_exc),
    .io_covSum(sfma_io_covSum),
    .metaAssert(sfma_metaAssert),
    .metaReset(sfma_metaReset),
    .fma_halt(sfma_fma_halt)
  );
  FPToInt fpiu ( // @[FPU.scala 763:20]
    .clock(fpiu_clock),
    .io_in_valid(fpiu_io_in_valid),
    .io_in_bits_ren2(fpiu_io_in_bits_ren2),
    .io_in_bits_singleIn(fpiu_io_in_bits_singleIn),
    .io_in_bits_singleOut(fpiu_io_in_bits_singleOut),
    .io_in_bits_wflags(fpiu_io_in_bits_wflags),
    .io_in_bits_rm(fpiu_io_in_bits_rm),
    .io_in_bits_typ(fpiu_io_in_bits_typ),
    .io_in_bits_in1(fpiu_io_in_bits_in1),
    .io_in_bits_in2(fpiu_io_in_bits_in2),
    .io_out_bits_in_rm(fpiu_io_out_bits_in_rm),
    .io_out_bits_in_in1(fpiu_io_out_bits_in_in1),
    .io_out_bits_in_in2(fpiu_io_out_bits_in_in2),
    .io_out_bits_lt(fpiu_io_out_bits_lt),
    .io_out_bits_store(fpiu_io_out_bits_store),
    .io_out_bits_toint(fpiu_io_out_bits_toint),
    .io_out_bits_exc(fpiu_io_out_bits_exc),
    .io_covSum(fpiu_io_covSum),
    .metaAssert(fpiu_metaAssert),
    .metaReset(fpiu_metaReset)
  );
  IntToFP ifpu ( // @[FPU.scala 773:20]
    .clock(ifpu_clock),
    .reset(ifpu_reset),
    .io_in_valid(ifpu_io_in_valid),
    .io_in_bits_singleIn(ifpu_io_in_bits_singleIn),
    .io_in_bits_wflags(ifpu_io_in_bits_wflags),
    .io_in_bits_rm(ifpu_io_in_bits_rm),
    .io_in_bits_typ(ifpu_io_in_bits_typ),
    .io_in_bits_in1(ifpu_io_in_bits_in1),
    .io_out_bits_data(ifpu_io_out_bits_data),
    .io_out_bits_exc(ifpu_io_out_bits_exc),
    .io_covSum(ifpu_io_covSum),
    .metaAssert(ifpu_metaAssert),
    .metaReset(ifpu_metaReset)
  );
  FPToFP fpmu ( // @[FPU.scala 778:20]
    .clock(fpmu_clock),
    .reset(fpmu_reset),
    .io_in_valid(fpmu_io_in_valid),
    .io_in_bits_ren2(fpmu_io_in_bits_ren2),
    .io_in_bits_singleOut(fpmu_io_in_bits_singleOut),
    .io_in_bits_wflags(fpmu_io_in_bits_wflags),
    .io_in_bits_rm(fpmu_io_in_bits_rm),
    .io_in_bits_in1(fpmu_io_in_bits_in1),
    .io_in_bits_in2(fpmu_io_in_bits_in2),
    .io_out_bits_data(fpmu_io_out_bits_data),
    .io_out_bits_exc(fpmu_io_out_bits_exc),
    .io_lt(fpmu_io_lt),
    .io_covSum(fpmu_io_covSum),
    .metaAssert(fpmu_metaAssert),
    .metaReset(fpmu_metaReset)
  );
  FPUFMAPipe_1 dfma ( // @[FPU.scala 797:28]
    .clock(dfma_clock),
    .reset(dfma_reset),
    .io_in_valid(dfma_io_in_valid),
    .io_in_bits_ren3(dfma_io_in_bits_ren3),
    .io_in_bits_swap23(dfma_io_in_bits_swap23),
    .io_in_bits_rm(dfma_io_in_bits_rm),
    .io_in_bits_fmaCmd(dfma_io_in_bits_fmaCmd),
    .io_in_bits_in1(dfma_io_in_bits_in1),
    .io_in_bits_in2(dfma_io_in_bits_in2),
    .io_in_bits_in3(dfma_io_in_bits_in3),
    .io_out_bits_data(dfma_io_out_bits_data),
    .io_out_bits_exc(dfma_io_out_bits_exc),
    .io_covSum(dfma_io_covSum),
    .metaAssert(dfma_metaAssert),
    .metaReset(dfma_metaReset),
    .fma_halt(dfma_fma_halt)
  );
  DivSqrtRecFN_small divSqrt ( // @[FPU.scala 887:27]
    .clock(divSqrt_clock),
    .reset(divSqrt_reset),
    .io_inReady(divSqrt_io_inReady),
    .io_inValid(divSqrt_io_inValid),
    .io_sqrtOp(divSqrt_io_sqrtOp),
    .io_a(divSqrt_io_a),
    .io_b(divSqrt_io_b),
    .io_roundingMode(divSqrt_io_roundingMode),
    .io_outValid_div(divSqrt_io_outValid_div),
    .io_outValid_sqrt(divSqrt_io_outValid_sqrt),
    .io_out(divSqrt_io_out),
    .io_exceptionFlags(divSqrt_io_exceptionFlags),
    .io_covSum(divSqrt_io_covSum),
    .metaAssert(divSqrt_metaAssert),
    .metaReset(divSqrt_metaReset),
    .divSqrtRecFNToRaw_halt(divSqrt_divSqrtRecFNToRaw_halt)
  );
  DivSqrtRecFN_small_1 divSqrt_1 ( // @[FPU.scala 887:27]
    .clock(divSqrt_1_clock),
    .reset(divSqrt_1_reset),
    .io_inReady(divSqrt_1_io_inReady),
    .io_inValid(divSqrt_1_io_inValid),
    .io_sqrtOp(divSqrt_1_io_sqrtOp),
    .io_a(divSqrt_1_io_a),
    .io_b(divSqrt_1_io_b),
    .io_roundingMode(divSqrt_1_io_roundingMode),
    .io_outValid_div(divSqrt_1_io_outValid_div),
    .io_outValid_sqrt(divSqrt_1_io_outValid_sqrt),
    .io_out(divSqrt_1_io_out),
    .io_exceptionFlags(divSqrt_1_io_exceptionFlags),
    .io_covSum(divSqrt_1_io_covSum),
    .metaAssert(divSqrt_1_metaAssert),
    .metaReset(divSqrt_1_metaReset),
    .divSqrtRecFNToRaw_halt(divSqrt_1_divSqrtRecFNToRaw_halt)
  );
  assign regfile__T_499_addr = ex_ra_0;
  assign regfile__T_499_data = regfile[regfile__T_499_addr]; // @[FPU.scala 715:20]
  assign regfile__T_502_addr = ex_ra_1;
  assign regfile__T_502_data = regfile[regfile__T_502_addr]; // @[FPU.scala 715:20]
  assign regfile__T_505_addr = ex_ra_2;
  assign regfile__T_505_data = regfile[regfile__T_505_addr]; // @[FPU.scala 715:20]
  assign regfile__T_472_data = _T_471 ? _T_468 : _T_311;
  assign regfile__T_472_addr = load_wb_tag;
  assign regfile__T_472_mask = 1'h1;
  assign regfile__T_472_en = load_wb;
  assign regfile__T_1002_data = wdouble ? _T_952 : _T_963;
  assign regfile__T_1002_addr = divSqrt_wen ? divSqrt_waddr : wbInfo_0_rd;
  assign regfile__T_1002_mask = 1'h1;
  assign regfile__T_1002_en = wen[0] | divSqrt_wen;
  assign killm = io_killm | io_nack_mem; // @[FPU.scala 690:25]
  assign _T_47 = mem_reg_valid & killm; // @[FPU.scala 694:41]
  assign killx = io_killx | _T_47; // @[FPU.scala 694:24]
  assign _T_49 = ex_reg_valid & ~killx; // @[FPU.scala 695:33]
  assign _T_54 = mem_reg_valid & ~killm; // @[FPU.scala 697:45]
  assign _T_67 = load_wb_double ? 64'h0 : 64'hffffffff00000000; // @[package.scala 31:71]
  assign _T_68 = _T_67 | load_wb_data; // @[FPU.scala 358:23]
  assign _T_72 = _T_68[62:52] == 11'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_73 = _T_68[51:0] == 52'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_78 = {{16'd0}, _T_68[31:16]}; // @[Bitwise.scala 103:31]
  assign _T_80 = {_T_68[15:0], 16'h0}; // @[Bitwise.scala 103:65]
  assign _T_82 = _T_80 & 32'hffff0000; // @[Bitwise.scala 103:75]
  assign _T_83 = _T_78 | _T_82; // @[Bitwise.scala 103:39]
  assign _GEN_165 = {{8'd0}, _T_83[31:8]}; // @[Bitwise.scala 103:31]
  assign _T_88 = _GEN_165 & 32'hff00ff; // @[Bitwise.scala 103:31]
  assign _T_90 = {_T_83[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_92 = _T_90 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  assign _T_93 = _T_88 | _T_92; // @[Bitwise.scala 103:39]
  assign _GEN_166 = {{4'd0}, _T_93[31:4]}; // @[Bitwise.scala 103:31]
  assign _T_98 = _GEN_166 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  assign _T_100 = {_T_93[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_102 = _T_100 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  assign _T_103 = _T_98 | _T_102; // @[Bitwise.scala 103:39]
  assign _GEN_167 = {{2'd0}, _T_103[31:2]}; // @[Bitwise.scala 103:31]
  assign _T_108 = _GEN_167 & 32'h33333333; // @[Bitwise.scala 103:31]
  assign _T_110 = {_T_103[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_112 = _T_110 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  assign _T_113 = _T_108 | _T_112; // @[Bitwise.scala 103:39]
  assign _GEN_168 = {{1'd0}, _T_113[31:1]}; // @[Bitwise.scala 103:31]
  assign _T_118 = _GEN_168 & 32'h55555555; // @[Bitwise.scala 103:31]
  assign _T_120 = {_T_113[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_122 = _T_120 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  assign _T_123 = _T_118 | _T_122; // @[Bitwise.scala 103:39]
  assign _T_129 = {{8'd0}, _T_68[47:40]}; // @[Bitwise.scala 103:31]
  assign _T_131 = {_T_68[39:32], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_133 = _T_131 & 16'hff00; // @[Bitwise.scala 103:75]
  assign _T_134 = _T_129 | _T_133; // @[Bitwise.scala 103:39]
  assign _GEN_169 = {{4'd0}, _T_134[15:4]}; // @[Bitwise.scala 103:31]
  assign _T_139 = _GEN_169 & 16'hf0f; // @[Bitwise.scala 103:31]
  assign _T_141 = {_T_134[11:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_143 = _T_141 & 16'hf0f0; // @[Bitwise.scala 103:75]
  assign _T_144 = _T_139 | _T_143; // @[Bitwise.scala 103:39]
  assign _GEN_170 = {{2'd0}, _T_144[15:2]}; // @[Bitwise.scala 103:31]
  assign _T_149 = _GEN_170 & 16'h3333; // @[Bitwise.scala 103:31]
  assign _T_151 = {_T_144[13:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_153 = _T_151 & 16'hcccc; // @[Bitwise.scala 103:75]
  assign _T_154 = _T_149 | _T_153; // @[Bitwise.scala 103:39]
  assign _GEN_171 = {{1'd0}, _T_154[15:1]}; // @[Bitwise.scala 103:31]
  assign _T_159 = _GEN_171 & 16'h5555; // @[Bitwise.scala 103:31]
  assign _T_161 = {_T_154[14:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_163 = _T_161 & 16'haaaa; // @[Bitwise.scala 103:75]
  assign _T_164 = _T_159 | _T_163; // @[Bitwise.scala 103:39]
  assign _T_176 = {_T_123,_T_164,_T_68[48],_T_68[49],_T_68[50],_T_68[51]}; // @[Cat.scala 30:58]
  assign _T_229 = _T_176[50] ? 6'h32 : 6'h33; // @[Mux.scala 31:69]
  assign _T_230 = _T_176[49] ? 6'h31 : _T_229; // @[Mux.scala 31:69]
  assign _T_231 = _T_176[48] ? 6'h30 : _T_230; // @[Mux.scala 31:69]
  assign _T_232 = _T_176[47] ? 6'h2f : _T_231; // @[Mux.scala 31:69]
  assign _T_233 = _T_176[46] ? 6'h2e : _T_232; // @[Mux.scala 31:69]
  assign _T_234 = _T_176[45] ? 6'h2d : _T_233; // @[Mux.scala 31:69]
  assign _T_235 = _T_176[44] ? 6'h2c : _T_234; // @[Mux.scala 31:69]
  assign _T_236 = _T_176[43] ? 6'h2b : _T_235; // @[Mux.scala 31:69]
  assign _T_237 = _T_176[42] ? 6'h2a : _T_236; // @[Mux.scala 31:69]
  assign _T_238 = _T_176[41] ? 6'h29 : _T_237; // @[Mux.scala 31:69]
  assign _T_239 = _T_176[40] ? 6'h28 : _T_238; // @[Mux.scala 31:69]
  assign _T_240 = _T_176[39] ? 6'h27 : _T_239; // @[Mux.scala 31:69]
  assign _T_241 = _T_176[38] ? 6'h26 : _T_240; // @[Mux.scala 31:69]
  assign _T_242 = _T_176[37] ? 6'h25 : _T_241; // @[Mux.scala 31:69]
  assign _T_243 = _T_176[36] ? 6'h24 : _T_242; // @[Mux.scala 31:69]
  assign _T_244 = _T_176[35] ? 6'h23 : _T_243; // @[Mux.scala 31:69]
  assign _T_245 = _T_176[34] ? 6'h22 : _T_244; // @[Mux.scala 31:69]
  assign _T_246 = _T_176[33] ? 6'h21 : _T_245; // @[Mux.scala 31:69]
  assign _T_247 = _T_176[32] ? 6'h20 : _T_246; // @[Mux.scala 31:69]
  assign _T_248 = _T_176[31] ? 6'h1f : _T_247; // @[Mux.scala 31:69]
  assign _T_249 = _T_176[30] ? 6'h1e : _T_248; // @[Mux.scala 31:69]
  assign _T_250 = _T_176[29] ? 6'h1d : _T_249; // @[Mux.scala 31:69]
  assign _T_251 = _T_176[28] ? 6'h1c : _T_250; // @[Mux.scala 31:69]
  assign _T_252 = _T_176[27] ? 6'h1b : _T_251; // @[Mux.scala 31:69]
  assign _T_253 = _T_176[26] ? 6'h1a : _T_252; // @[Mux.scala 31:69]
  assign _T_254 = _T_176[25] ? 6'h19 : _T_253; // @[Mux.scala 31:69]
  assign _T_255 = _T_176[24] ? 6'h18 : _T_254; // @[Mux.scala 31:69]
  assign _T_256 = _T_176[23] ? 6'h17 : _T_255; // @[Mux.scala 31:69]
  assign _T_257 = _T_176[22] ? 6'h16 : _T_256; // @[Mux.scala 31:69]
  assign _T_258 = _T_176[21] ? 6'h15 : _T_257; // @[Mux.scala 31:69]
  assign _T_259 = _T_176[20] ? 6'h14 : _T_258; // @[Mux.scala 31:69]
  assign _T_260 = _T_176[19] ? 6'h13 : _T_259; // @[Mux.scala 31:69]
  assign _T_261 = _T_176[18] ? 6'h12 : _T_260; // @[Mux.scala 31:69]
  assign _T_262 = _T_176[17] ? 6'h11 : _T_261; // @[Mux.scala 31:69]
  assign _T_263 = _T_176[16] ? 6'h10 : _T_262; // @[Mux.scala 31:69]
  assign _T_264 = _T_176[15] ? 6'hf : _T_263; // @[Mux.scala 31:69]
  assign _T_265 = _T_176[14] ? 6'he : _T_264; // @[Mux.scala 31:69]
  assign _T_266 = _T_176[13] ? 6'hd : _T_265; // @[Mux.scala 31:69]
  assign _T_267 = _T_176[12] ? 6'hc : _T_266; // @[Mux.scala 31:69]
  assign _T_268 = _T_176[11] ? 6'hb : _T_267; // @[Mux.scala 31:69]
  assign _T_269 = _T_176[10] ? 6'ha : _T_268; // @[Mux.scala 31:69]
  assign _T_270 = _T_176[9] ? 6'h9 : _T_269; // @[Mux.scala 31:69]
  assign _T_271 = _T_176[8] ? 6'h8 : _T_270; // @[Mux.scala 31:69]
  assign _T_272 = _T_176[7] ? 6'h7 : _T_271; // @[Mux.scala 31:69]
  assign _T_273 = _T_176[6] ? 6'h6 : _T_272; // @[Mux.scala 31:69]
  assign _T_274 = _T_176[5] ? 6'h5 : _T_273; // @[Mux.scala 31:69]
  assign _T_275 = _T_176[4] ? 6'h4 : _T_274; // @[Mux.scala 31:69]
  assign _T_276 = _T_176[3] ? 6'h3 : _T_275; // @[Mux.scala 31:69]
  assign _T_277 = _T_176[2] ? 6'h2 : _T_276; // @[Mux.scala 31:69]
  assign _T_278 = _T_176[1] ? 6'h1 : _T_277; // @[Mux.scala 31:69]
  assign _T_279 = _T_176[0] ? 6'h0 : _T_278; // @[Mux.scala 31:69]
  assign _GEN_172 = {{63'd0}, _T_68[51:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_280 = _GEN_172 << _T_279; // @[rawFloatFromFN.scala 54:36]
  assign _T_282 = {_T_280[50:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_173 = {{6'd0}, _T_279}; // @[rawFloatFromFN.scala 57:26]
  assign _T_283 = _GEN_173 ^ 12'hfff; // @[rawFloatFromFN.scala 57:26]
  assign _T_284 = _T_72 ? _T_283 : {{1'd0}, _T_68[62:52]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_285 = _T_72 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_174 = {{9'd0}, _T_285}; // @[rawFloatFromFN.scala 60:22]
  assign _T_286 = 11'h400 | _GEN_174; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_175 = {{1'd0}, _T_286}; // @[rawFloatFromFN.scala 59:15]
  assign _T_288 = _T_284 + _GEN_175; // @[rawFloatFromFN.scala 59:15]
  assign _T_289 = _T_72 & _T_73; // @[rawFloatFromFN.scala 62:34]
  assign _T_291 = _T_288[11:10] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_295 = _T_291 & ~_T_73; // @[rawFloatFromFN.scala 66:33]
  assign _T_298 = {1'b0,$signed(_T_288)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_300 = _T_72 ? _T_282 : _T_68[51:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_302 = {1'h0,~_T_289,_T_300}; // @[Cat.scala 30:58]
  assign _T_304 = _T_289 ? 3'h0 : _T_298[11:9]; // @[recFNFromFN.scala 48:16]
  assign _GEN_176 = {{2'd0}, _T_295}; // @[recFNFromFN.scala 48:79]
  assign _T_306 = _T_304 | _GEN_176; // @[recFNFromFN.scala 48:79]
  assign _T_311 = {_T_68[63],_T_306,_T_298[8:0],_T_302[51:0]}; // @[Cat.scala 30:58]
  assign _T_315 = _T_68[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_316 = _T_68[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_321 = {{8'd0}, _T_68[15:8]}; // @[Bitwise.scala 103:31]
  assign _T_323 = {_T_68[7:0], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_325 = _T_323 & 16'hff00; // @[Bitwise.scala 103:75]
  assign _T_326 = _T_321 | _T_325; // @[Bitwise.scala 103:39]
  assign _GEN_177 = {{4'd0}, _T_326[15:4]}; // @[Bitwise.scala 103:31]
  assign _T_331 = _GEN_177 & 16'hf0f; // @[Bitwise.scala 103:31]
  assign _T_333 = {_T_326[11:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_335 = _T_333 & 16'hf0f0; // @[Bitwise.scala 103:75]
  assign _T_336 = _T_331 | _T_335; // @[Bitwise.scala 103:39]
  assign _GEN_178 = {{2'd0}, _T_336[15:2]}; // @[Bitwise.scala 103:31]
  assign _T_341 = _GEN_178 & 16'h3333; // @[Bitwise.scala 103:31]
  assign _T_343 = {_T_336[13:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_345 = _T_343 & 16'hcccc; // @[Bitwise.scala 103:75]
  assign _T_346 = _T_341 | _T_345; // @[Bitwise.scala 103:39]
  assign _GEN_179 = {{1'd0}, _T_346[15:1]}; // @[Bitwise.scala 103:31]
  assign _T_351 = _GEN_179 & 16'h5555; // @[Bitwise.scala 103:31]
  assign _T_353 = {_T_346[14:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_355 = _T_353 & 16'haaaa; // @[Bitwise.scala 103:75]
  assign _T_356 = _T_351 | _T_355; // @[Bitwise.scala 103:39]
  assign _T_376 = {_T_356,_T_68[16],_T_68[17],_T_68[18],_T_68[19],_T_68[20],_T_68[21],_T_68[22]}; // @[Cat.scala 30:58]
  assign _T_400 = _T_376[21] ? 5'h15 : 5'h16; // @[Mux.scala 31:69]
  assign _T_401 = _T_376[20] ? 5'h14 : _T_400; // @[Mux.scala 31:69]
  assign _T_402 = _T_376[19] ? 5'h13 : _T_401; // @[Mux.scala 31:69]
  assign _T_403 = _T_376[18] ? 5'h12 : _T_402; // @[Mux.scala 31:69]
  assign _T_404 = _T_376[17] ? 5'h11 : _T_403; // @[Mux.scala 31:69]
  assign _T_405 = _T_376[16] ? 5'h10 : _T_404; // @[Mux.scala 31:69]
  assign _T_406 = _T_376[15] ? 5'hf : _T_405; // @[Mux.scala 31:69]
  assign _T_407 = _T_376[14] ? 5'he : _T_406; // @[Mux.scala 31:69]
  assign _T_408 = _T_376[13] ? 5'hd : _T_407; // @[Mux.scala 31:69]
  assign _T_409 = _T_376[12] ? 5'hc : _T_408; // @[Mux.scala 31:69]
  assign _T_410 = _T_376[11] ? 5'hb : _T_409; // @[Mux.scala 31:69]
  assign _T_411 = _T_376[10] ? 5'ha : _T_410; // @[Mux.scala 31:69]
  assign _T_412 = _T_376[9] ? 5'h9 : _T_411; // @[Mux.scala 31:69]
  assign _T_413 = _T_376[8] ? 5'h8 : _T_412; // @[Mux.scala 31:69]
  assign _T_414 = _T_376[7] ? 5'h7 : _T_413; // @[Mux.scala 31:69]
  assign _T_415 = _T_376[6] ? 5'h6 : _T_414; // @[Mux.scala 31:69]
  assign _T_416 = _T_376[5] ? 5'h5 : _T_415; // @[Mux.scala 31:69]
  assign _T_417 = _T_376[4] ? 5'h4 : _T_416; // @[Mux.scala 31:69]
  assign _T_418 = _T_376[3] ? 5'h3 : _T_417; // @[Mux.scala 31:69]
  assign _T_419 = _T_376[2] ? 5'h2 : _T_418; // @[Mux.scala 31:69]
  assign _T_420 = _T_376[1] ? 5'h1 : _T_419; // @[Mux.scala 31:69]
  assign _T_421 = _T_376[0] ? 5'h0 : _T_420; // @[Mux.scala 31:69]
  assign _GEN_180 = {{31'd0}, _T_68[22:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_422 = _GEN_180 << _T_421; // @[rawFloatFromFN.scala 54:36]
  assign _T_424 = {_T_422[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_181 = {{4'd0}, _T_421}; // @[rawFloatFromFN.scala 57:26]
  assign _T_425 = _GEN_181 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  assign _T_426 = _T_315 ? _T_425 : {{1'd0}, _T_68[30:23]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_427 = _T_315 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_182 = {{6'd0}, _T_427}; // @[rawFloatFromFN.scala 60:22]
  assign _T_428 = 8'h80 | _GEN_182; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_183 = {{1'd0}, _T_428}; // @[rawFloatFromFN.scala 59:15]
  assign _T_430 = _T_426 + _GEN_183; // @[rawFloatFromFN.scala 59:15]
  assign _T_431 = _T_315 & _T_316; // @[rawFloatFromFN.scala 62:34]
  assign _T_433 = _T_430[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_437 = _T_433 & ~_T_316; // @[rawFloatFromFN.scala 66:33]
  assign _T_440 = {1'b0,$signed(_T_430)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_442 = _T_315 ? _T_424 : _T_68[22:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_444 = {1'h0,~_T_431,_T_442}; // @[Cat.scala 30:58]
  assign _T_446 = _T_431 ? 3'h0 : _T_440[8:6]; // @[recFNFromFN.scala 48:16]
  assign _GEN_184 = {{2'd0}, _T_437}; // @[recFNFromFN.scala 48:79]
  assign _T_448 = _T_446 | _GEN_184; // @[recFNFromFN.scala 48:79]
  assign _T_453 = {_T_68[31],_T_448,_T_440[5:0],_T_444[22:0]}; // @[Cat.scala 30:58]
  assign _T_457 = ~_T_311[51:32] == 20'h0; // @[FPU.scala 265:42]
  assign _T_468 = {_T_311[64:61],_T_457,_T_311[59:53],_T_453[31],_T_311[51:32],_T_453[32],_T_453[30:0]}; // @[Cat.scala 30:58]
  assign _T_471 = ~_T_311[63:61] == 3'h0; // @[FPU.scala 197:56]
  assign wdata = _T_471 ? _T_468 : _T_311; // @[FPU.scala 271:8]
  assign _T_485 = ~wdata[63:61] == 3'h0; // @[FPU.scala 197:56]
  assign _T_490 = ~wdata[51:32] == 20'h0; // @[FPU.scala 312:96]
  assign _T_491 = wdata[60] == _T_490; // @[FPU.scala 312:55]
  assign _T_492 = ~_T_485 | _T_491; // @[FPU.scala 312:31]
  assign _T_495 = _T_492 | reset; // @[FPU.scala 719:11]
  assign _T_513 = ~fp_decoder_io_sigs_swap12 & ~fp_decoder_io_sigs_swap23; // @[FPU.scala 733:29]
  assign _T_517 = ex_reg_inst[14:12] == 3'h7; // @[FPU.scala 737:38]
  assign _T_519 = ex_reg_valid & ex_reg_ctrl_fma; // @[FPU.scala 760:33]
  assign tag = ~ex_reg_ctrl_singleIn; // @[FPU.scala 741:15]
  assign _T_526 = {regfile__T_499_data[31],regfile__T_499_data[52],regfile__T_499_data[30:0]}; // @[Cat.scala 30:58]
  assign _T_529 = ~regfile__T_499_data[64:60] == 5'h0; // @[FPU.scala 259:84]
  assign _T_551 = _T_529 ? 33'h0 : 33'he0400000; // @[FPU.scala 299:31]
  assign _T_552 = _T_526 | _T_551; // @[FPU.scala 299:26]
  assign _T_557 = {regfile__T_502_data[31],regfile__T_502_data[52],regfile__T_502_data[30:0]}; // @[Cat.scala 30:58]
  assign _T_560 = ~regfile__T_502_data[64:60] == 5'h0; // @[FPU.scala 259:84]
  assign _T_582 = _T_560 ? 33'h0 : 33'he0400000; // @[FPU.scala 299:31]
  assign _T_583 = _T_557 | _T_582; // @[FPU.scala 299:26]
  assign _T_588 = {regfile__T_505_data[31],regfile__T_505_data[52],regfile__T_505_data[30:0]}; // @[Cat.scala 30:58]
  assign _T_591 = ~regfile__T_505_data[64:60] == 5'h0; // @[FPU.scala 259:84]
  assign _T_613 = _T_591 ? 33'h0 : 33'he0400000; // @[FPU.scala 299:31]
  assign _T_614 = _T_588 | _T_613; // @[FPU.scala 299:26]
  assign _T_619 = ~ex_reg_ctrl_ren3 & ex_reg_inst[27]; // @[FPU.scala 748:53]
  assign _GEN_185 = {{1'd0}, _T_619}; // @[FPU.scala 748:36]
  assign _T_621 = ex_reg_ctrl_toint | ex_reg_ctrl_div; // @[FPU.scala 764:51]
  assign _T_622 = _T_621 | ex_reg_ctrl_sqrt; // @[FPU.scala 764:66]
  assign _T_623 = ex_reg_ctrl_fastpipe & ex_reg_ctrl_wflags; // @[FPU.scala 764:103]
  assign _T_624 = _T_622 | _T_623; // @[FPU.scala 764:82]
  assign _T_635 = {_T_526[22:0], 53'h0}; // @[FPU.scala 225:28]
  assign _GEN_186 = {{3'd0}, _T_526[31:23]}; // @[FPU.scala 228:31]
  assign _T_639 = _GEN_186 + 12'h800; // @[FPU.scala 228:31]
  assign _T_642 = _T_639 - 12'h100; // @[FPU.scala 228:48]
  assign _T_643 = _T_526[31:29] == 3'h0; // @[FPU.scala 229:19]
  assign _T_644 = _T_526[31:29] >= 3'h6; // @[FPU.scala 229:36]
  assign _T_645 = _T_643 | _T_644; // @[FPU.scala 229:25]
  assign _T_647 = {_T_526[31:29],_T_642[8:0]}; // @[Cat.scala 30:58]
  assign _T_649 = _T_645 ? _T_647 : _T_642; // @[FPU.scala 229:10]
  assign _T_651 = {_T_526[32],_T_649,_T_635[75:24]}; // @[Cat.scala 30:58]
  assign _T_657 = tag | _T_529; // @[package.scala 31:71]
  assign _T_659 = tag ? regfile__T_499_data : _T_651; // @[package.scala 31:71]
  assign _T_669 = {_T_557[22:0], 53'h0}; // @[FPU.scala 225:28]
  assign _GEN_187 = {{3'd0}, _T_557[31:23]}; // @[FPU.scala 228:31]
  assign _T_673 = _GEN_187 + 12'h800; // @[FPU.scala 228:31]
  assign _T_676 = _T_673 - 12'h100; // @[FPU.scala 228:48]
  assign _T_677 = _T_557[31:29] == 3'h0; // @[FPU.scala 229:19]
  assign _T_678 = _T_557[31:29] >= 3'h6; // @[FPU.scala 229:36]
  assign _T_679 = _T_677 | _T_678; // @[FPU.scala 229:25]
  assign _T_681 = {_T_557[31:29],_T_676[8:0]}; // @[Cat.scala 30:58]
  assign _T_683 = _T_679 ? _T_681 : _T_676; // @[FPU.scala 229:10]
  assign _T_685 = {_T_557[32],_T_683,_T_669[75:24]}; // @[Cat.scala 30:58]
  assign _T_691 = tag | _T_560; // @[package.scala 31:71]
  assign _T_693 = tag ? regfile__T_502_data : _T_685; // @[package.scala 31:71]
  assign _T_738 = {{1'd0}, io_fromint_data}; // @[FPU.scala 776:29]
  assign _T_851 = mem_ctrl_fma & mem_ctrl_singleOut; // @[FPU.scala 795:56]
  assign _T_852 = _T_851 ? 2'h2 : 2'h0; // @[FPU.scala 804:23]
  assign _T_854 = mem_ctrl_fma & ~mem_ctrl_singleOut; // @[FPU.scala 800:62]
  assign _T_855 = _T_854 ? 3'h4 : 3'h0; // @[FPU.scala 804:23]
  assign _T_856 = mem_ctrl_fastpipe | mem_ctrl_fromint; // @[FPU.scala 804:78]
  assign _GEN_194 = {{1'd0}, _T_856}; // @[FPU.scala 804:78]
  assign _T_857 = _GEN_194 | _T_852; // @[FPU.scala 804:78]
  assign _GEN_195 = {{1'd0}, _T_857}; // @[FPU.scala 804:78]
  assign memLatencyMask = _GEN_195 | _T_855; // @[FPU.scala 804:78]
  assign _T_867 = mem_ctrl_fma | mem_ctrl_fastpipe; // @[FPU.scala 820:48]
  assign _T_868 = _T_867 | mem_ctrl_fromint; // @[FPU.scala 820:69]
  assign mem_wen = mem_reg_valid & _T_868; // @[FPU.scala 820:31]
  assign _T_869 = ex_reg_ctrl_fastpipe ? 2'h2 : 2'h0; // @[FPU.scala 804:23]
  assign _T_870 = ex_reg_ctrl_fromint ? 2'h2 : 2'h0; // @[FPU.scala 804:23]
  assign _T_871 = ex_reg_ctrl_fma & ex_reg_ctrl_singleOut; // @[FPU.scala 795:56]
  assign _T_872 = _T_871 ? 3'h4 : 3'h0; // @[FPU.scala 804:23]
  assign _T_874 = ex_reg_ctrl_fma & ~ex_reg_ctrl_singleOut; // @[FPU.scala 800:62]
  assign _T_875 = _T_874 ? 4'h8 : 4'h0; // @[FPU.scala 804:23]
  assign _T_876 = _T_869 | _T_870; // @[FPU.scala 804:78]
  assign _GEN_196 = {{1'd0}, _T_876}; // @[FPU.scala 804:78]
  assign _T_877 = _GEN_196 | _T_872; // @[FPU.scala 804:78]
  assign _GEN_197 = {{1'd0}, _T_877}; // @[FPU.scala 804:78]
  assign _T_878 = _GEN_197 | _T_875; // @[FPU.scala 804:78]
  assign _GEN_198 = {{1'd0}, memLatencyMask}; // @[FPU.scala 821:62]
  assign _T_879 = _GEN_198 & _T_878; // @[FPU.scala 821:62]
  assign _T_880 = _T_879 != 4'h0; // @[FPU.scala 821:89]
  assign _T_881 = mem_wen & _T_880; // @[FPU.scala 821:43]
  assign _T_882 = ex_reg_ctrl_fastpipe ? 3'h4 : 3'h0; // @[FPU.scala 804:23]
  assign _T_883 = ex_reg_ctrl_fromint ? 3'h4 : 3'h0; // @[FPU.scala 804:23]
  assign _T_885 = _T_871 ? 4'h8 : 4'h0; // @[FPU.scala 804:23]
  assign _T_888 = _T_874 ? 5'h10 : 5'h0; // @[FPU.scala 804:23]
  assign _T_889 = _T_882 | _T_883; // @[FPU.scala 804:78]
  assign _GEN_199 = {{1'd0}, _T_889}; // @[FPU.scala 804:78]
  assign _T_890 = _GEN_199 | _T_885; // @[FPU.scala 804:78]
  assign _GEN_200 = {{1'd0}, _T_890}; // @[FPU.scala 804:78]
  assign _T_891 = _GEN_200 | _T_888; // @[FPU.scala 804:78]
  assign _GEN_201 = {{2'd0}, wen}; // @[FPU.scala 821:101]
  assign _T_892 = _GEN_201 & _T_891; // @[FPU.scala 821:101]
  assign _T_893 = _T_892 != 5'h0; // @[FPU.scala 821:128]
  assign _T_894 = _T_881 | _T_893; // @[FPU.scala 821:93]
  assign _GEN_202 = {{1'd0}, wen[2:1]}; // @[FPU.scala 830:23]
  assign _T_902 = _GEN_202 | memLatencyMask; // @[FPU.scala 830:23]
  assign _T_905 = ~write_port_busy & memLatencyMask[0]; // @[FPU.scala 833:30]
  assign _T_912 = _T_854 ? 2'h3 : 2'h0; // @[FPU.scala 806:63]
  assign _GEN_203 = {{1'd0}, mem_ctrl_fromint}; // @[FPU.scala 806:108]
  assign _T_914 = _GEN_203 | _T_852; // @[FPU.scala 806:108]
  assign _T_915 = _T_914 | _T_912; // @[FPU.scala 806:108]
  assign _T_919 = ~write_port_busy & memLatencyMask[1]; // @[FPU.scala 833:30]
  assign _T_933 = ~write_port_busy & memLatencyMask[2]; // @[FPU.scala 833:30]
  assign divSqrt_typeTag = divSqrt_1_io_outValid_div | divSqrt_1_io_outValid_sqrt; // @[FPU.scala 902:37]
  assign _T_1111 = divSqrt_io_outValid_div | divSqrt_io_outValid_sqrt; // @[FPU.scala 902:37]
  assign _GEN_154 = _T_1111 & ~divSqrt_killed; // @[FPU.scala 902:66]
  assign divSqrt_wen = divSqrt_typeTag ? ~divSqrt_killed : _GEN_154; // @[FPU.scala 902:66]
  assign wdouble = divSqrt_wen ? divSqrt_typeTag : ~wbInfo_0_single; // @[FPU.scala 843:20]
  assign _T_946 = wbInfo_0_pipeid == 2'h1; // @[package.scala 31:81]
  assign _T_947 = _T_946 ? ifpu_io_out_bits_data : fpmu_io_out_bits_data; // @[package.scala 31:71]
  assign _T_948 = wbInfo_0_pipeid == 2'h2; // @[package.scala 31:81]
  assign _T_949 = _T_948 ? sfma_io_out_bits_data : _T_947; // @[package.scala 31:71]
  assign _T_950 = wbInfo_0_pipeid == 2'h3; // @[package.scala 31:81]
  assign _T_951 = _T_950 ? dfma_io_out_bits_data : _T_949; // @[package.scala 31:71]
  assign _T_1128 = ~divSqrt_1_io_out[63:61] == 3'h0; // @[FPU.scala 197:56]
  assign _T_1125 = divSqrt_1_io_out & 65'h1efefffffffffffff; // @[FPU.scala 340:25]
  assign _T_1129 = _T_1128 ? _T_1125 : divSqrt_1_io_out; // @[FPU.scala 341:10]
  assign _GEN_155 = divSqrt_io_out; // @[FPU.scala 902:66]
  assign divSqrt_wdata = divSqrt_typeTag ? _T_1129 : {{32'd0}, _GEN_155}; // @[FPU.scala 902:66]
  assign _T_952 = divSqrt_wen ? divSqrt_wdata : _T_951; // @[FPU.scala 844:22]
  assign _T_963 = {5'h1f,7'h7f,_T_952[31],20'hfffff,_T_952[32],_T_952[30:0]}; // @[Cat.scala 30:58]
  assign wdata_1 = wdouble ? _T_952 : _T_963; // @[package.scala 31:71]
  assign _T_970 = _T_946 ? ifpu_io_out_bits_exc : fpmu_io_out_bits_exc; // @[package.scala 31:71]
  assign _T_972 = _T_948 ? sfma_io_out_bits_exc : _T_970; // @[package.scala 31:71]
  assign wexc = _T_950 ? dfma_io_out_bits_exc : _T_972; // @[package.scala 31:71]
  assign _T_977 = wen[0] | divSqrt_wen; // @[FPU.scala 846:35]
  assign _T_990 = ~wdata_1[63:61] == 3'h0; // @[FPU.scala 197:56]
  assign _T_995 = ~wdata_1[51:32] == 20'h0; // @[FPU.scala 312:96]
  assign _T_996 = wdata_1[60] == _T_995; // @[FPU.scala 312:55]
  assign _T_997 = ~_T_990 | _T_996; // @[FPU.scala 312:31]
  assign _T_1000 = _T_997 | reset; // @[FPU.scala 847:11]
  assign wb_toint_valid = wb_reg_valid & wb_ctrl_toint; // @[FPU.scala 859:37]
  assign _T_1007 = wb_toint_valid | divSqrt_wen; // @[FPU.scala 861:41]
  assign _T_1010 = wb_toint_valid ? wb_toint_exc : 5'h0; // @[FPU.scala 863:8]
  assign _GEN_156 = divSqrt_io_exceptionFlags; // @[FPU.scala 902:66]
  assign divSqrt_flags = divSqrt_typeTag ? divSqrt_1_io_exceptionFlags : _GEN_156; // @[FPU.scala 902:66]
  assign _T_1011 = divSqrt_wen ? divSqrt_flags : 5'h0; // @[FPU.scala 864:8]
  assign _T_1012 = _T_1010 | _T_1011; // @[FPU.scala 863:48]
  assign _T_1014 = wen[0] ? wexc : 5'h0; // @[FPU.scala 865:8]
  assign _T_1016 = mem_ctrl_div | mem_ctrl_sqrt; // @[FPU.scala 867:47]
  assign _T_1017 = wen != 3'h0; // @[FPU.scala 867:72]
  assign divSqrt_write_port_busy = _T_1016 & _T_1017; // @[FPU.scala 867:65]
  assign _T_1018 = ex_reg_valid & ex_reg_ctrl_wflags; // @[FPU.scala 868:33]
  assign _T_1019 = mem_reg_valid & mem_ctrl_wflags; // @[FPU.scala 868:68]
  assign _T_1020 = _T_1018 | _T_1019; // @[FPU.scala 868:51]
  assign _T_1022 = _T_1020 | wb_toint_valid; // @[FPU.scala 868:87]
  assign _T_1024 = _T_1022 | _T_1017; // @[FPU.scala 868:120]
  assign divSqrt_inFlight = ~divSqrt_1_io_inReady | ~divSqrt_io_inReady; // @[FPU.scala 895:34]
  assign _T_1025 = _T_1024 | divSqrt_inFlight; // @[FPU.scala 868:131]
  assign _T_1027 = write_port_busy | divSqrt_write_port_busy; // @[FPU.scala 869:34]
  assign _T_1034 = _T_854 | mem_ctrl_div; // @[FPU.scala 872:96]
  assign _T_1043 = wen[0] & _T_950; // @[FPU.scala 873:60]
  assign _T_1048 = io_inst[14:12] == 3'h5; // @[package.scala 14:47]
  assign _T_1049 = io_inst[14:12] == 3'h6; // @[package.scala 14:47]
  assign _T_1050 = _T_1048 | _T_1049; // @[package.scala 14:62]
  assign _T_1052 = io_inst[14:12] == 3'h7; // @[FPU.scala 877:67]
  assign _T_1053 = io_fcsr_rm >= 3'h5; // @[FPU.scala 877:87]
  assign _T_1054 = _T_1052 & _T_1053; // @[FPU.scala 877:73]
  assign _T_1063 = mem_reg_valid & mem_ctrl_singleOut; // @[FPU.scala 888:43]
  assign _T_1065 = _T_1063 & _T_1016; // @[FPU.scala 888:65]
  assign _T_1071 = {fpiu_io_out_bits_in_in1[51:0], 24'h0}; // @[FPU.scala 225:28]
  assign _T_1075 = fpiu_io_out_bits_in_in1[63:52] + 12'h100; // @[FPU.scala 228:31]
  assign _T_1078 = _T_1075 - 12'h800; // @[FPU.scala 228:48]
  assign _T_1079 = fpiu_io_out_bits_in_in1[63:61] == 3'h0; // @[FPU.scala 229:19]
  assign _T_1080 = fpiu_io_out_bits_in_in1[63:61] >= 3'h6; // @[FPU.scala 229:36]
  assign _T_1081 = _T_1079 | _T_1080; // @[FPU.scala 229:25]
  assign _T_1083 = {fpiu_io_out_bits_in_in1[63:61],_T_1078[5:0]}; // @[Cat.scala 30:58]
  assign _T_1085 = _T_1081 ? _T_1083 : _T_1078[8:0]; // @[FPU.scala 229:10]
  assign _T_1086 = {fpiu_io_out_bits_in_in1[64],_T_1085}; // @[Cat.scala 30:58]
  assign _T_1091 = {fpiu_io_out_bits_in_in2[51:0], 24'h0}; // @[FPU.scala 225:28]
  assign _T_1095 = fpiu_io_out_bits_in_in2[63:52] + 12'h100; // @[FPU.scala 228:31]
  assign _T_1098 = _T_1095 - 12'h800; // @[FPU.scala 228:48]
  assign _T_1099 = fpiu_io_out_bits_in_in2[63:61] == 3'h0; // @[FPU.scala 229:19]
  assign _T_1100 = fpiu_io_out_bits_in_in2[63:61] >= 3'h6; // @[FPU.scala 229:36]
  assign _T_1101 = _T_1099 | _T_1100; // @[FPU.scala 229:25]
  assign _T_1103 = {fpiu_io_out_bits_in_in2[63:61],_T_1098[5:0]}; // @[Cat.scala 30:58]
  assign _T_1105 = _T_1101 ? _T_1103 : _T_1098[8:0]; // @[FPU.scala 229:10]
  assign _T_1106 = {fpiu_io_out_bits_in_in2[64],_T_1105}; // @[Cat.scala 30:58]
  assign _T_1109 = divSqrt_io_inValid & divSqrt_io_inReady; // @[FPU.scala 897:32]
  assign _T_1114 = mem_reg_valid & ~mem_ctrl_singleOut; // @[FPU.scala 888:43]
  assign _T_1116 = _T_1114 & _T_1016; // @[FPU.scala 888:65]
  assign _T_1120 = divSqrt_1_io_inValid & divSqrt_1_io_inReady; // @[FPU.scala 897:32]
  assign io_fcsr_flags_valid = _T_1007 | wen[0]; // @[FPU.scala 861:23]
  assign io_fcsr_flags_bits = _T_1012 | _T_1014; // @[FPU.scala 862:22]
  assign io_store_data = fpiu_io_out_bits_store; // @[FPU.scala 766:17]
  assign io_toint_data = fpiu_io_out_bits_toint; // @[FPU.scala 767:17]
  assign io_fcsr_rdy = ~_T_1025; // @[FPU.scala 868:15]
  assign io_nack_mem = _T_1027 | divSqrt_inFlight; // @[FPU.scala 869:15]
  assign io_illegal_rm = _T_1050 | _T_1054; // @[FPU.scala 877:17]
  assign io_dec_wen = fp_decoder_io_sigs_wen; // @[FPU.scala 870:10]
  assign io_dec_ren1 = fp_decoder_io_sigs_ren1; // @[FPU.scala 870:10]
  assign io_dec_ren2 = fp_decoder_io_sigs_ren2; // @[FPU.scala 870:10]
  assign io_dec_ren3 = fp_decoder_io_sigs_ren3; // @[FPU.scala 870:10]
  assign io_sboard_set = wb_reg_valid & _T_1037; // @[FPU.scala 872:17]
  assign io_sboard_clr = divSqrt_wen | _T_1043; // @[FPU.scala 873:17]
  assign io_sboard_clra = divSqrt_wen ? divSqrt_waddr : wbInfo_0_rd; // @[FPU.scala 874:18]
  assign fp_decoder_io_inst = io_inst; // @[FPU.scala 675:22]
  assign sfma_clock = clock;
  assign sfma_reset = reset;
  assign sfma_io_in_valid = _T_519 & ex_reg_ctrl_singleOut; // @[FPU.scala 760:20]
  assign sfma_io_in_bits_ren3 = ex_reg_ctrl_ren3; // @[FPU.scala 761:19]
  assign sfma_io_in_bits_swap23 = ex_reg_ctrl_swap23; // @[FPU.scala 761:19]
  assign sfma_io_in_bits_rm = _T_517 ? io_fcsr_rm : ex_reg_inst[14:12]; // @[FPU.scala 761:19]
  assign sfma_io_in_bits_fmaCmd = ex_reg_inst[3:2] | _GEN_185; // @[FPU.scala 761:19]
  assign sfma_io_in_bits_in1 = {{32'd0}, _T_552}; // @[FPU.scala 761:19]
  assign sfma_io_in_bits_in2 = {{32'd0}, _T_583}; // @[FPU.scala 761:19]
  assign sfma_io_in_bits_in3 = {{32'd0}, _T_614}; // @[FPU.scala 761:19]
  assign fpiu_clock = clock;
  assign fpiu_io_in_valid = ex_reg_valid & _T_624; // @[FPU.scala 764:20]
  assign fpiu_io_in_bits_ren2 = ex_reg_ctrl_ren2; // @[FPU.scala 765:19]
  assign fpiu_io_in_bits_singleIn = ex_reg_ctrl_singleIn; // @[FPU.scala 765:19]
  assign fpiu_io_in_bits_singleOut = ex_reg_ctrl_singleOut; // @[FPU.scala 765:19]
  assign fpiu_io_in_bits_wflags = ex_reg_ctrl_wflags; // @[FPU.scala 765:19]
  assign fpiu_io_in_bits_rm = _T_517 ? io_fcsr_rm : ex_reg_inst[14:12]; // @[FPU.scala 765:19]
  assign fpiu_io_in_bits_typ = ex_reg_inst[21:20]; // @[FPU.scala 765:19]
  assign fpiu_io_in_bits_in1 = _T_657 ? _T_659 : 65'he008000000000000; // @[FPU.scala 765:19]
  assign fpiu_io_in_bits_in2 = _T_691 ? _T_693 : 65'he008000000000000; // @[FPU.scala 765:19]
  assign ifpu_clock = clock;
  assign ifpu_reset = reset;
  assign ifpu_io_in_valid = ex_reg_valid & ex_reg_ctrl_fromint; // @[FPU.scala 774:20]
  assign ifpu_io_in_bits_singleIn = fpiu_io_in_bits_singleIn; // @[FPU.scala 775:19]
  assign ifpu_io_in_bits_wflags = fpiu_io_in_bits_wflags; // @[FPU.scala 775:19]
  assign ifpu_io_in_bits_rm = fpiu_io_in_bits_rm; // @[FPU.scala 775:19]
  assign ifpu_io_in_bits_typ = fpiu_io_in_bits_typ; // @[FPU.scala 775:19]
  assign ifpu_io_in_bits_in1 = _T_738[63:0]; // @[FPU.scala 775:19 FPU.scala 776:23]
  assign fpmu_clock = clock;
  assign fpmu_reset = reset;
  assign fpmu_io_in_valid = ex_reg_valid & ex_reg_ctrl_fastpipe; // @[FPU.scala 779:20]
  assign fpmu_io_in_bits_ren2 = fpiu_io_in_bits_ren2; // @[FPU.scala 780:19]
  assign fpmu_io_in_bits_singleOut = fpiu_io_in_bits_singleOut; // @[FPU.scala 780:19]
  assign fpmu_io_in_bits_wflags = fpiu_io_in_bits_wflags; // @[FPU.scala 780:19]
  assign fpmu_io_in_bits_rm = fpiu_io_in_bits_rm; // @[FPU.scala 780:19]
  assign fpmu_io_in_bits_in1 = fpiu_io_in_bits_in1; // @[FPU.scala 780:19]
  assign fpmu_io_in_bits_in2 = fpiu_io_in_bits_in2; // @[FPU.scala 780:19]
  assign fpmu_io_lt = fpiu_io_out_bits_lt; // @[FPU.scala 781:14]
  assign dfma_clock = clock;
  assign dfma_reset = reset;
  assign dfma_io_in_valid = _T_519 & ~ex_reg_ctrl_singleOut; // @[FPU.scala 798:28]
  assign dfma_io_in_bits_ren3 = ex_reg_ctrl_ren3; // @[FPU.scala 799:27]
  assign dfma_io_in_bits_swap23 = ex_reg_ctrl_swap23; // @[FPU.scala 799:27]
  assign dfma_io_in_bits_rm = _T_517 ? io_fcsr_rm : ex_reg_inst[14:12]; // @[FPU.scala 799:27]
  assign dfma_io_in_bits_fmaCmd = ex_reg_inst[3:2] | _GEN_185; // @[FPU.scala 799:27]
  assign dfma_io_in_bits_in1 = regfile__T_499_data; // @[FPU.scala 799:27]
  assign dfma_io_in_bits_in2 = regfile__T_502_data; // @[FPU.scala 799:27]
  assign dfma_io_in_bits_in3 = regfile__T_505_data; // @[FPU.scala 799:27]
  assign divSqrt_clock = clock;
  assign divSqrt_reset = reset;
  assign divSqrt_io_inValid = _T_1065 & ~divSqrt_inFlight; // @[FPU.scala 888:26]
  assign divSqrt_io_sqrtOp = mem_ctrl_sqrt; // @[FPU.scala 889:25]
  assign divSqrt_io_a = {_T_1086,_T_1071[75:53]}; // @[FPU.scala 890:20]
  assign divSqrt_io_b = {_T_1106,_T_1091[75:53]}; // @[FPU.scala 891:20]
  assign divSqrt_io_roundingMode = fpiu_io_out_bits_in_rm; // @[FPU.scala 892:31]
  assign divSqrt_1_clock = clock;
  assign divSqrt_1_reset = reset;
  assign divSqrt_1_io_inValid = _T_1116 & ~divSqrt_inFlight; // @[FPU.scala 888:26]
  assign divSqrt_1_io_sqrtOp = mem_ctrl_sqrt; // @[FPU.scala 889:25]
  assign divSqrt_1_io_a = fpiu_io_out_bits_in_in1; // @[FPU.scala 890:20]
  assign divSqrt_1_io_b = fpiu_io_out_bits_in_in2; // @[FPU.scala 891:20]
  assign divSqrt_1_io_roundingMode = fpiu_io_out_bits_in_rm; // @[FPU.scala 892:31]
  assign FPU_cov_read_addr = FPU_state;
  assign FPU_cov_read_data = FPU_cov[FPU_cov_read_addr]; // @[Coverage map for FPU]
  assign FPU_cov_write_data = 1'h1;
  assign FPU_cov_write_addr = FPU_state;
  assign FPU_cov_write_mask = 1'h1;
  assign FPU_cov_write_en = 1'h1;
  assign wen_shl = {wen, 14'h0};
  assign wen_pad = {3'h0,wen_shl};
  assign wb_reg_valid_shl = {wb_reg_valid, 16'h0};
  assign wb_reg_valid_pad = {3'h0,wb_reg_valid_shl};
  assign ex_reg_valid_shl = {ex_reg_valid, 18'h0};
  assign ex_reg_valid_pad = {1'h0,ex_reg_valid_shl};
  assign mem_ctrl_fma_shl = {mem_ctrl_fma, 7'h0};
  assign mem_ctrl_fma_pad = {12'h0,mem_ctrl_fma_shl};
  assign mem_ctrl_fromint_shl = {mem_ctrl_fromint, 14'h0};
  assign mem_ctrl_fromint_pad = {5'h0,mem_ctrl_fromint_shl};
  assign wbInfo_0_pipeid_shl = {wbInfo_0_pipeid, 15'h0};
  assign wbInfo_0_pipeid_pad = {3'h0,wbInfo_0_pipeid_shl};
  assign ex_reg_ctrl_fma_shl = {ex_reg_ctrl_fma, 3'h0};
  assign ex_reg_ctrl_fma_pad = {16'h0,ex_reg_ctrl_fma_shl};
  assign mem_reg_valid_shl = {mem_reg_valid, 19'h0};
  assign mem_reg_valid_pad = mem_reg_valid_shl;
  assign ex_reg_ctrl_singleIn_shl = {ex_reg_ctrl_singleIn, 15'h0};
  assign ex_reg_ctrl_singleIn_pad = {4'h0,ex_reg_ctrl_singleIn_shl};
  assign wbInfo_0_single_shl = {wbInfo_0_single, 1'h0};
  assign wbInfo_0_single_pad = {18'h0,wbInfo_0_single_shl};
  assign mem_ctrl_singleOut_shl = {mem_ctrl_singleOut, 14'h0};
  assign mem_ctrl_singleOut_pad = {5'h0,mem_ctrl_singleOut_shl};
  assign ex_reg_ctrl_singleOut_shl = {ex_reg_ctrl_singleOut, 11'h0};
  assign ex_reg_ctrl_singleOut_pad = {8'h0,ex_reg_ctrl_singleOut_shl};
  assign mem_ctrl_toint_shl = {mem_ctrl_toint, 18'h0};
  assign mem_ctrl_toint_pad = {1'h0,mem_ctrl_toint_shl};
  assign ex_reg_ctrl_fromint_shl = {ex_reg_ctrl_fromint, 6'h0};
  assign ex_reg_ctrl_fromint_pad = {13'h0,ex_reg_ctrl_fromint_shl};
  assign ex_reg_ctrl_fastpipe_shl = {ex_reg_ctrl_fastpipe, 8'h0};
  assign ex_reg_ctrl_fastpipe_pad = {11'h0,ex_reg_ctrl_fastpipe_shl};
  assign mem_ctrl_fastpipe_shl = {mem_ctrl_fastpipe, 6'h0};
  assign mem_ctrl_fastpipe_pad = {13'h0,mem_ctrl_fastpipe_shl};
  assign write_port_busy_shl = {write_port_busy, 9'h0};
  assign write_port_busy_pad = {10'h0,write_port_busy_shl};
  assign load_wb_double_shl = {load_wb_double, 4'h0};
  assign load_wb_double_pad = {15'h0,load_wb_double_shl};
  assign divSqrt_killed_shl = {divSqrt_killed, 10'h0};
  assign divSqrt_killed_pad = {9'h0,divSqrt_killed_shl};
  assign wb_ctrl_toint_shl = {wb_ctrl_toint, 2'h0};
  assign wb_ctrl_toint_pad = {17'h0,wb_ctrl_toint_shl};
  assign FPU_xor7 = wen_pad ^ wb_reg_valid_pad;
  assign FPU_xor18 = mem_ctrl_fma_pad ^ mem_ctrl_fromint_pad;
  assign FPU_xor8 = ex_reg_valid_pad ^ FPU_xor18;
  assign FPU_xor3 = FPU_xor7 ^ FPU_xor8;
  assign FPU_xor9 = wbInfo_0_pipeid_pad ^ ex_reg_ctrl_fma_pad;
  assign FPU_xor22 = ex_reg_ctrl_singleIn_pad ^ wbInfo_0_single_pad;
  assign FPU_xor10 = mem_reg_valid_pad ^ FPU_xor22;
  assign FPU_xor4 = FPU_xor9 ^ FPU_xor10;
  assign FPU_xor1 = FPU_xor3 ^ FPU_xor4;
  assign FPU_xor11 = mem_ctrl_singleOut_pad ^ ex_reg_ctrl_singleOut_pad;
  assign FPU_xor26 = ex_reg_ctrl_fromint_pad ^ ex_reg_ctrl_fastpipe_pad;
  assign FPU_xor12 = mem_ctrl_toint_pad ^ FPU_xor26;
  assign FPU_xor5 = FPU_xor11 ^ FPU_xor12;
  assign FPU_xor13 = mem_ctrl_fastpipe_pad ^ write_port_busy_pad;
  assign FPU_xor30 = divSqrt_killed_pad ^ wb_ctrl_toint_pad;
  assign FPU_xor14 = load_wb_double_pad ^ FPU_xor30;
  assign FPU_xor6 = FPU_xor13 ^ FPU_xor14;
  assign FPU_xor2 = FPU_xor5 ^ FPU_xor6;
  assign FPU_xor0 = FPU_xor1 ^ FPU_xor2;
  assign fp_decoder_sum = FPU_covSum + fp_decoder_io_covSum;
  assign dfma_sum = fp_decoder_sum + dfma_io_covSum;
  assign fpmu_sum = dfma_sum + fpmu_io_covSum;
  assign divSqrt_1_sum = fpmu_sum + divSqrt_1_io_covSum;
  assign ifpu_sum = divSqrt_1_sum + ifpu_io_covSum;
  assign divSqrt_sum = ifpu_sum + divSqrt_io_covSum;
  assign fpiu_sum = divSqrt_sum + fpiu_io_covSum;
  assign sfma_sum = fpiu_sum + sfma_io_covSum;
  assign io_covSum = sfma_sum;
  assign stopEn0 = load_wb & ~_T_495;
  assign stopEn1 = _T_977 & ~_T_1000;
  assign divSqrt_metaAssert_wire = divSqrt_metaAssert;
  assign dfma_metaAssert_wire = dfma_metaAssert;
  assign fpiu_metaAssert_wire = fpiu_metaAssert;
  assign fpmu_metaAssert_wire = fpmu_metaAssert;
  assign divSqrt_1_metaAssert_wire = divSqrt_1_metaAssert;
  assign sfma_metaAssert_wire = sfma_metaAssert;
  assign ifpu_metaAssert_wire = ifpu_metaAssert;
  assign fp_decoder_metaAssert_wire = fp_decoder_metaAssert;
  assign FPU_or3 = stopEn0 | stopEn1;
  assign FPU_or10 = divSqrt_metaAssert_wire | divSqrt_1_metaAssert_wire;
  assign FPU_or4 = fp_decoder_metaAssert_wire | FPU_or10;
  assign FPU_or1 = FPU_or3 | FPU_or4;
  assign FPU_or5 = fpiu_metaAssert_wire | dfma_metaAssert_wire;
  assign FPU_or14 = ifpu_metaAssert_wire | sfma_metaAssert_wire;
  assign FPU_or6 = fpmu_metaAssert_wire | FPU_or14;
  assign FPU_or2 = FPU_or5 | FPU_or6;
  assign FPU_or0 = FPU_or1 | FPU_or2;
  assign metaAssert = FPU_metaAssert;
  assign dfma_metaReset = metaReset | dfma_halt;
  assign fpmu_metaReset = metaReset | fpmu_halt;
  assign divSqrt_1_metaReset = metaReset | divSqrt_1_halt;
  assign ifpu_metaReset = metaReset | ifpu_halt;
  assign divSqrt_metaReset = metaReset | divSqrt_halt;
  assign fpiu_metaReset = metaReset | fpiu_halt;
  assign sfma_metaReset = metaReset | sfma_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {3{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regfile[initvar] = _RAND_0[64:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ex_reg_valid = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ex_reg_inst = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ex_reg_ctrl_ren2 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  ex_reg_ctrl_ren3 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  ex_reg_ctrl_swap23 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  ex_reg_ctrl_singleIn = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ex_reg_ctrl_singleOut = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  ex_reg_ctrl_fromint = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  ex_reg_ctrl_toint = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  ex_reg_ctrl_fastpipe = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  ex_reg_ctrl_fma = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  ex_reg_ctrl_div = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  ex_reg_ctrl_sqrt = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  ex_reg_ctrl_wflags = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  ex_ra_0 = _RAND_15[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  ex_ra_1 = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  ex_ra_2 = _RAND_17[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  mem_reg_valid = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  mem_reg_inst = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  wb_reg_valid = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  mem_ctrl_singleOut = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  mem_ctrl_fromint = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  mem_ctrl_toint = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  mem_ctrl_fastpipe = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  mem_ctrl_fma = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  mem_ctrl_div = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  mem_ctrl_sqrt = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  mem_ctrl_wflags = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  wb_ctrl_toint = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  load_wb = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  load_wb_double = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {2{`RANDOM}};
  load_wb_data = _RAND_32[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  load_wb_tag = _RAND_33[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  divSqrt_waddr = _RAND_34[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  wen = _RAND_35[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  wbInfo_0_rd = _RAND_36[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  wbInfo_0_single = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  wbInfo_0_pipeid = _RAND_38[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  wbInfo_1_rd = _RAND_39[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  wbInfo_1_single = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  wbInfo_1_pipeid = _RAND_41[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  wbInfo_2_rd = _RAND_42[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  wbInfo_2_single = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  wbInfo_2_pipeid = _RAND_44[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  write_port_busy = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  divSqrt_killed = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  wb_toint_exc = _RAND_47[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_1037 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  FPU_state = _RAND_49[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    FPU_cov[initvar] = _RAND_50[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  FPU_covSum = _RAND_51[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  FPU_metaAssert = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(regfile__T_472_en & regfile__T_472_mask) begin
      regfile[regfile__T_472_addr] <= regfile__T_472_data; // @[FPU.scala 715:20]
    end
    if(regfile__T_1002_en & regfile__T_1002_mask) begin
      regfile[regfile__T_1002_addr] <= regfile__T_1002_data; // @[FPU.scala 715:20]
    end
    if (metaReset) begin
      ex_reg_valid <= 1'h0;
    end else if (reset) begin
      ex_reg_valid <= 1'h0;
    end else begin
      ex_reg_valid <= io_valid;
    end
    if (metaReset) begin
      ex_reg_inst <= 32'h0;
    end else if (io_valid) begin
      ex_reg_inst <= io_inst;
    end
    if (metaReset) begin
      ex_reg_ctrl_ren2 <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_ren2 <= fp_decoder_io_sigs_ren2;
    end
    if (metaReset) begin
      ex_reg_ctrl_ren3 <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_ren3 <= fp_decoder_io_sigs_ren3;
    end
    if (metaReset) begin
      ex_reg_ctrl_swap23 <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_swap23 <= fp_decoder_io_sigs_swap23;
    end
    if (metaReset) begin
      ex_reg_ctrl_singleIn <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_singleIn <= fp_decoder_io_sigs_singleIn;
    end
    if (metaReset) begin
      ex_reg_ctrl_singleOut <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_singleOut <= fp_decoder_io_sigs_singleOut;
    end
    if (metaReset) begin
      ex_reg_ctrl_fromint <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_fromint <= fp_decoder_io_sigs_fromint;
    end
    if (metaReset) begin
      ex_reg_ctrl_toint <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_toint <= fp_decoder_io_sigs_toint;
    end
    if (metaReset) begin
      ex_reg_ctrl_fastpipe <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_fastpipe <= fp_decoder_io_sigs_fastpipe;
    end
    if (metaReset) begin
      ex_reg_ctrl_fma <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_fma <= fp_decoder_io_sigs_fma;
    end
    if (metaReset) begin
      ex_reg_ctrl_div <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_div <= fp_decoder_io_sigs_div;
    end
    if (metaReset) begin
      ex_reg_ctrl_sqrt <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_sqrt <= fp_decoder_io_sigs_sqrt;
    end
    if (metaReset) begin
      ex_reg_ctrl_wflags <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_wflags <= fp_decoder_io_sigs_wflags;
    end
    if (metaReset) begin
      ex_ra_0 <= 5'h0;
    end else if (io_valid) begin
      if (fp_decoder_io_sigs_ren2) begin
        if (fp_decoder_io_sigs_swap12) begin
          ex_ra_0 <= io_inst[24:20];
        end else if (fp_decoder_io_sigs_ren1) begin
          if (~fp_decoder_io_sigs_swap12) begin
            ex_ra_0 <= io_inst[19:15];
          end
        end
      end else if (fp_decoder_io_sigs_ren1) begin
        if (~fp_decoder_io_sigs_swap12) begin
          ex_ra_0 <= io_inst[19:15];
        end
      end
    end
    if (metaReset) begin
      ex_ra_1 <= 5'h0;
    end else if (io_valid) begin
      if (fp_decoder_io_sigs_ren2) begin
        if (_T_513) begin
          ex_ra_1 <= io_inst[24:20];
        end else if (fp_decoder_io_sigs_ren1) begin
          if (fp_decoder_io_sigs_swap12) begin
            ex_ra_1 <= io_inst[19:15];
          end
        end
      end else if (fp_decoder_io_sigs_ren1) begin
        if (fp_decoder_io_sigs_swap12) begin
          ex_ra_1 <= io_inst[19:15];
        end
      end
    end
    if (metaReset) begin
      ex_ra_2 <= 5'h0;
    end else if (io_valid) begin
      if (fp_decoder_io_sigs_ren3) begin
        ex_ra_2 <= io_inst[31:27];
      end else if (fp_decoder_io_sigs_ren2) begin
        if (fp_decoder_io_sigs_swap23) begin
          ex_ra_2 <= io_inst[24:20];
        end
      end
    end
    if (metaReset) begin
      mem_reg_valid <= 1'h0;
    end else if (reset) begin
      mem_reg_valid <= 1'h0;
    end else begin
      mem_reg_valid <= _T_49;
    end
    if (metaReset) begin
      mem_reg_inst <= 32'h0;
    end else if (ex_reg_valid) begin
      mem_reg_inst <= ex_reg_inst;
    end
    if (metaReset) begin
      wb_reg_valid <= 1'h0;
    end else if (reset) begin
      wb_reg_valid <= 1'h0;
    end else begin
      wb_reg_valid <= _T_54;
    end
    if (metaReset) begin
      mem_ctrl_singleOut <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_singleOut <= ex_reg_ctrl_singleOut;
    end
    if (metaReset) begin
      mem_ctrl_fromint <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_fromint <= ex_reg_ctrl_fromint;
    end
    if (metaReset) begin
      mem_ctrl_toint <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_toint <= ex_reg_ctrl_toint;
    end
    if (metaReset) begin
      mem_ctrl_fastpipe <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_fastpipe <= ex_reg_ctrl_fastpipe;
    end
    if (metaReset) begin
      mem_ctrl_fma <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_fma <= ex_reg_ctrl_fma;
    end
    if (metaReset) begin
      mem_ctrl_div <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_div <= ex_reg_ctrl_div;
    end
    if (metaReset) begin
      mem_ctrl_sqrt <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_sqrt <= ex_reg_ctrl_sqrt;
    end
    if (metaReset) begin
      mem_ctrl_wflags <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_wflags <= ex_reg_ctrl_wflags;
    end
    if (metaReset) begin
      wb_ctrl_toint <= 1'h0;
    end else if (mem_reg_valid) begin
      wb_ctrl_toint <= mem_ctrl_toint;
    end
    if (metaReset) begin
      load_wb <= 1'h0;
    end else begin
      load_wb <= io_dmem_resp_val;
    end
    if (metaReset) begin
      load_wb_double <= 1'h0;
    end else if (io_dmem_resp_val) begin
      load_wb_double <= io_dmem_resp_type[0];
    end
    if (metaReset) begin
      load_wb_data <= 64'h0;
    end else if (io_dmem_resp_val) begin
      load_wb_data <= io_dmem_resp_data;
    end
    if (metaReset) begin
      load_wb_tag <= 5'h0;
    end else if (io_dmem_resp_val) begin
      load_wb_tag <= io_dmem_resp_tag;
    end
    if (metaReset) begin
      divSqrt_waddr <= 5'h0;
    end else if (_T_1120) begin
      divSqrt_waddr <= mem_reg_inst[11:7];
    end else if (_T_1109) begin
      divSqrt_waddr <= mem_reg_inst[11:7];
    end
    if (metaReset) begin
      wen <= 3'h0;
    end else if (reset) begin
      wen <= 3'h0;
    end else if (mem_wen) begin
      if (~killm) begin
        wen <= _T_902;
      end else begin
        wen <= {{1'd0}, wen[2:1]};
      end
    end else begin
      wen <= {{1'd0}, wen[2:1]};
    end
    if (metaReset) begin
      wbInfo_0_rd <= 5'h0;
    end else if (mem_wen) begin
      if (_T_905) begin
        wbInfo_0_rd <= mem_reg_inst[11:7];
      end else if (wen[1]) begin
        wbInfo_0_rd <= wbInfo_1_rd;
      end
    end else if (wen[1]) begin
      wbInfo_0_rd <= wbInfo_1_rd;
    end
    if (metaReset) begin
      wbInfo_0_single <= 1'h0;
    end else if (mem_wen) begin
      if (_T_905) begin
        wbInfo_0_single <= mem_ctrl_singleOut;
      end else if (wen[1]) begin
        wbInfo_0_single <= wbInfo_1_single;
      end
    end else if (wen[1]) begin
      wbInfo_0_single <= wbInfo_1_single;
    end
    if (metaReset) begin
      wbInfo_0_pipeid <= 2'h0;
    end else if (mem_wen) begin
      if (_T_905) begin
        wbInfo_0_pipeid <= _T_915;
      end else if (wen[1]) begin
        wbInfo_0_pipeid <= wbInfo_1_pipeid;
      end
    end else if (wen[1]) begin
      wbInfo_0_pipeid <= wbInfo_1_pipeid;
    end
    if (metaReset) begin
      wbInfo_1_rd <= 5'h0;
    end else if (mem_wen) begin
      if (_T_919) begin
        wbInfo_1_rd <= mem_reg_inst[11:7];
      end else if (wen[2]) begin
        wbInfo_1_rd <= wbInfo_2_rd;
      end
    end else if (wen[2]) begin
      wbInfo_1_rd <= wbInfo_2_rd;
    end
    if (metaReset) begin
      wbInfo_1_single <= 1'h0;
    end else if (mem_wen) begin
      if (_T_919) begin
        wbInfo_1_single <= mem_ctrl_singleOut;
      end else if (wen[2]) begin
        wbInfo_1_single <= wbInfo_2_single;
      end
    end else if (wen[2]) begin
      wbInfo_1_single <= wbInfo_2_single;
    end
    if (metaReset) begin
      wbInfo_1_pipeid <= 2'h0;
    end else if (mem_wen) begin
      if (_T_919) begin
        wbInfo_1_pipeid <= _T_915;
      end else if (wen[2]) begin
        wbInfo_1_pipeid <= wbInfo_2_pipeid;
      end
    end else if (wen[2]) begin
      wbInfo_1_pipeid <= wbInfo_2_pipeid;
    end
    if (metaReset) begin
      wbInfo_2_rd <= 5'h0;
    end else if (mem_wen) begin
      if (_T_933) begin
        wbInfo_2_rd <= mem_reg_inst[11:7];
      end
    end
    if (metaReset) begin
      wbInfo_2_single <= 1'h0;
    end else if (mem_wen) begin
      if (_T_933) begin
        wbInfo_2_single <= mem_ctrl_singleOut;
      end
    end
    if (metaReset) begin
      wbInfo_2_pipeid <= 2'h0;
    end else if (mem_wen) begin
      if (_T_933) begin
        wbInfo_2_pipeid <= _T_915;
      end
    end
    if (metaReset) begin
      write_port_busy <= 1'h0;
    end else if (ex_reg_valid) begin
      write_port_busy <= _T_894;
    end
    if (metaReset) begin
      divSqrt_killed <= 1'h0;
    end else if (_T_1120) begin
      divSqrt_killed <= killm;
    end else if (_T_1109) begin
      divSqrt_killed <= killm;
    end
    if (metaReset) begin
      wb_toint_exc <= 5'h0;
    end else if (mem_ctrl_toint) begin
      wb_toint_exc <= fpiu_io_out_bits_exc;
    end
    if (metaReset) begin
      _T_1037 <= 1'h0;
    end else begin
      _T_1037 <= _T_1034 | mem_ctrl_sqrt;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (load_wb & ~_T_495) begin
          $fwrite(32'h80000002,"Assertion failed\n    at FPU.scala:719 assert(consistent(wdata))\n"); // @[FPU.scala 719:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (load_wb & ~_T_495) begin
          $fatal; // @[FPU.scala 719:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_977 & ~_T_1000) begin
          $fwrite(32'h80000002,"Assertion failed\n    at FPU.scala:847 assert(consistent(wdata))\n"); // @[FPU.scala 847:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_977 & ~_T_1000) begin
          $fatal; // @[FPU.scala 847:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    FPU_state <= FPU_xor0;
    if (!(FPU_cov_read_data)) begin
      FPU_covSum <= FPU_covSum + 1'h1;
    end
    if (metaReset) begin
      FPU_metaAssert <= 1'h0;
    end else begin
      FPU_metaAssert <= FPU_metaAssert | FPU_or0;
    end
  end
  always @(posedge clock) begin
    if(FPU_cov_write_en & FPU_cov_write_mask) begin
      FPU_cov[FPU_cov_write_addr] <= FPU_cov_write_data; // @[Coverage map for FPU]
    end
  end
endmodule
module HellaCacheArbiter(
  input         clock,
  output        io_requestor_0_req_ready,
  input         io_requestor_0_req_valid,
  input  [39:0] io_requestor_0_req_bits_addr,
  input         io_requestor_0_s1_kill,
  output        io_requestor_0_s2_nack,
  output        io_requestor_0_resp_valid,
  output [63:0] io_requestor_0_resp_bits_data_word_bypass,
  output        io_requestor_0_s2_xcpt_ae_ld,
  output        io_requestor_1_req_ready,
  input         io_requestor_1_req_valid,
  input  [39:0] io_requestor_1_req_bits_addr,
  input  [6:0]  io_requestor_1_req_bits_tag,
  input  [4:0]  io_requestor_1_req_bits_cmd,
  input  [2:0]  io_requestor_1_req_bits_typ,
  input         io_requestor_1_s1_kill,
  input  [63:0] io_requestor_1_s1_data_data,
  output        io_requestor_1_s2_nack,
  output        io_requestor_1_resp_valid,
  output [6:0]  io_requestor_1_resp_bits_tag,
  output [2:0]  io_requestor_1_resp_bits_typ,
  output [63:0] io_requestor_1_resp_bits_data,
  output        io_requestor_1_resp_bits_replay,
  output        io_requestor_1_resp_bits_has_data,
  output [63:0] io_requestor_1_resp_bits_data_word_bypass,
  output        io_requestor_1_replay_next,
  output        io_requestor_1_s2_xcpt_ma_ld,
  output        io_requestor_1_s2_xcpt_ma_st,
  output        io_requestor_1_s2_xcpt_pf_ld,
  output        io_requestor_1_s2_xcpt_pf_st,
  output        io_requestor_1_s2_xcpt_ae_ld,
  output        io_requestor_1_s2_xcpt_ae_st,
  output        io_requestor_1_ordered,
  output        io_requestor_1_perf_grant,
  input         io_requestor_1_keep_clock_enabled,
  output        io_requestor_1_clock_enabled,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [39:0] io_mem_req_bits_addr,
  output [6:0]  io_mem_req_bits_tag,
  output [4:0]  io_mem_req_bits_cmd,
  output [2:0]  io_mem_req_bits_typ,
  output        io_mem_req_bits_phys,
  output        io_mem_s1_kill,
  output [63:0] io_mem_s1_data_data,
  input         io_mem_s2_nack,
  input         io_mem_resp_valid,
  input  [6:0]  io_mem_resp_bits_tag,
  input  [2:0]  io_mem_resp_bits_typ,
  input  [63:0] io_mem_resp_bits_data,
  input         io_mem_resp_bits_replay,
  input         io_mem_resp_bits_has_data,
  input  [63:0] io_mem_resp_bits_data_word_bypass,
  input         io_mem_replay_next,
  input         io_mem_s2_xcpt_ma_ld,
  input         io_mem_s2_xcpt_ma_st,
  input         io_mem_s2_xcpt_pf_ld,
  input         io_mem_s2_xcpt_pf_st,
  input         io_mem_s2_xcpt_ae_ld,
  input         io_mem_s2_xcpt_ae_st,
  input         io_mem_ordered,
  input         io_mem_perf_grant,
  output        io_mem_keep_clock_enabled,
  input         io_mem_clock_enabled,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg  _T_210; // @[HellaCacheArbiter.scala 19:20]
  reg [31:0] _RAND_0;
  reg  _T_212; // @[HellaCacheArbiter.scala 20:20]
  reg [31:0] _RAND_1;
  wire [7:0] _T_217; // @[Cat.scala 30:58]
  wire [7:0] _GEN_4; // @[HellaCacheArbiter.scala 52:26]
  reg  HellaCacheArbiter_state; // @[Register tracking HellaCacheArbiter state]
  reg [31:0] _RAND_2;
  reg  HellaCacheArbiter_cov [0:1]; // @[Coverage map for HellaCacheArbiter]
  reg [31:0] _RAND_3;
  wire  HellaCacheArbiter_cov_read_data; // @[Coverage map for HellaCacheArbiter]
  wire  HellaCacheArbiter_cov_read_addr; // @[Coverage map for HellaCacheArbiter]
  wire  HellaCacheArbiter_cov_write_data; // @[Coverage map for HellaCacheArbiter]
  wire  HellaCacheArbiter_cov_write_addr; // @[Coverage map for HellaCacheArbiter]
  wire  HellaCacheArbiter_cov_write_mask; // @[Coverage map for HellaCacheArbiter]
  wire  HellaCacheArbiter_cov_write_en; // @[Coverage map for HellaCacheArbiter]
  reg [29:0] HellaCacheArbiter_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_4;
  wire  _T_210_shl;
  wire  _T_210_pad;
  assign _T_217 = {io_requestor_1_req_bits_tag,1'h1}; // @[Cat.scala 30:58]
  assign _GEN_4 = io_requestor_0_req_valid ? 8'h0 : _T_217; // @[HellaCacheArbiter.scala 52:26]
  assign io_requestor_0_req_ready = io_mem_req_ready; // @[HellaCacheArbiter.scala 25:31]
  assign io_requestor_0_s2_nack = io_mem_s2_nack & ~_T_212; // @[HellaCacheArbiter.scala 65:31]
  assign io_requestor_0_resp_valid = io_mem_resp_valid & ~io_mem_resp_bits_tag[0]; // @[HellaCacheArbiter.scala 61:18]
  assign io_requestor_0_resp_bits_data_word_bypass = io_mem_resp_bits_data_word_bypass; // @[HellaCacheArbiter.scala 68:17]
  assign io_requestor_0_s2_xcpt_ae_ld = io_mem_s2_xcpt_ae_ld; // @[HellaCacheArbiter.scala 62:31]
  assign io_requestor_1_req_ready = io_requestor_0_req_ready & ~io_requestor_0_req_valid; // @[HellaCacheArbiter.scala 27:33]
  assign io_requestor_1_s2_nack = io_mem_s2_nack & _T_212; // @[HellaCacheArbiter.scala 65:31]
  assign io_requestor_1_resp_valid = io_mem_resp_valid & io_mem_resp_bits_tag[0]; // @[HellaCacheArbiter.scala 61:18]
  assign io_requestor_1_resp_bits_tag = {{1'd0}, io_mem_resp_bits_tag[6:1]}; // @[HellaCacheArbiter.scala 68:17 HellaCacheArbiter.scala 69:21]
  assign io_requestor_1_resp_bits_typ = io_mem_resp_bits_typ; // @[HellaCacheArbiter.scala 68:17]
  assign io_requestor_1_resp_bits_data = io_mem_resp_bits_data; // @[HellaCacheArbiter.scala 68:17]
  assign io_requestor_1_resp_bits_replay = io_mem_resp_bits_replay; // @[HellaCacheArbiter.scala 68:17]
  assign io_requestor_1_resp_bits_has_data = io_mem_resp_bits_has_data; // @[HellaCacheArbiter.scala 68:17]
  assign io_requestor_1_resp_bits_data_word_bypass = io_mem_resp_bits_data_word_bypass; // @[HellaCacheArbiter.scala 68:17]
  assign io_requestor_1_replay_next = io_mem_replay_next; // @[HellaCacheArbiter.scala 71:35]
  assign io_requestor_1_s2_xcpt_ma_ld = io_mem_s2_xcpt_ma_ld; // @[HellaCacheArbiter.scala 62:31]
  assign io_requestor_1_s2_xcpt_ma_st = io_mem_s2_xcpt_ma_st; // @[HellaCacheArbiter.scala 62:31]
  assign io_requestor_1_s2_xcpt_pf_ld = io_mem_s2_xcpt_pf_ld; // @[HellaCacheArbiter.scala 62:31]
  assign io_requestor_1_s2_xcpt_pf_st = io_mem_s2_xcpt_pf_st; // @[HellaCacheArbiter.scala 62:31]
  assign io_requestor_1_s2_xcpt_ae_ld = io_mem_s2_xcpt_ae_ld; // @[HellaCacheArbiter.scala 62:31]
  assign io_requestor_1_s2_xcpt_ae_st = io_mem_s2_xcpt_ae_st; // @[HellaCacheArbiter.scala 62:31]
  assign io_requestor_1_ordered = io_mem_ordered; // @[HellaCacheArbiter.scala 63:31]
  assign io_requestor_1_perf_grant = io_mem_perf_grant; // @[HellaCacheArbiter.scala 64:28]
  assign io_requestor_1_clock_enabled = io_mem_clock_enabled; // @[HellaCacheArbiter.scala 67:37]
  assign io_mem_req_valid = io_requestor_0_req_valid | io_requestor_1_req_valid; // @[HellaCacheArbiter.scala 24:22]
  assign io_mem_req_bits_addr = io_requestor_0_req_valid ? io_requestor_0_req_bits_addr : io_requestor_1_req_bits_addr; // @[HellaCacheArbiter.scala 34:30 HellaCacheArbiter.scala 34:30]
  assign io_mem_req_bits_tag = _GEN_4[6:0]; // @[HellaCacheArbiter.scala 36:29 HellaCacheArbiter.scala 36:29]
  assign io_mem_req_bits_cmd = io_requestor_0_req_valid ? 5'h0 : io_requestor_1_req_bits_cmd; // @[HellaCacheArbiter.scala 32:29 HellaCacheArbiter.scala 32:29]
  assign io_mem_req_bits_typ = io_requestor_0_req_valid ? 3'h3 : io_requestor_1_req_bits_typ; // @[HellaCacheArbiter.scala 33:29 HellaCacheArbiter.scala 33:29]
  assign io_mem_req_bits_phys = io_requestor_0_req_valid; // @[HellaCacheArbiter.scala 35:30 HellaCacheArbiter.scala 35:30]
  assign io_mem_s1_kill = _T_210 ? io_requestor_1_s1_kill : io_requestor_0_s1_kill; // @[HellaCacheArbiter.scala 40:24 HellaCacheArbiter.scala 40:24]
  assign io_mem_s1_data_data = _T_210 ? io_requestor_1_s1_data_data : 64'h0; // @[HellaCacheArbiter.scala 41:24 HellaCacheArbiter.scala 41:24]
  assign io_mem_keep_clock_enabled = io_requestor_1_keep_clock_enabled; // @[HellaCacheArbiter.scala 22:31]
  assign HellaCacheArbiter_cov_read_addr = HellaCacheArbiter_state;
  assign HellaCacheArbiter_cov_read_data = HellaCacheArbiter_cov[HellaCacheArbiter_cov_read_addr]; // @[Coverage map for HellaCacheArbiter]
  assign HellaCacheArbiter_cov_write_data = 1'h1;
  assign HellaCacheArbiter_cov_write_addr = HellaCacheArbiter_state;
  assign HellaCacheArbiter_cov_write_mask = 1'h1;
  assign HellaCacheArbiter_cov_write_en = 1'h1;
  assign _T_210_shl = _T_210;
  assign _T_210_pad = _T_210_shl;
  assign io_covSum = HellaCacheArbiter_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_210 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_212 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  HellaCacheArbiter_state = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    HellaCacheArbiter_cov[initvar] = _RAND_3[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  HellaCacheArbiter_covSum = _RAND_4[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      _T_210 <= 1'h0;
    end else if (io_requestor_0_req_valid) begin
      _T_210 <= 1'h0;
    end else begin
      _T_210 <= 1'h1;
    end
    if (metaReset) begin
      _T_212 <= 1'h0;
    end else begin
      _T_212 <= _T_210;
    end
    HellaCacheArbiter_state <= _T_210_pad;
    if (!(HellaCacheArbiter_cov_read_data)) begin
      HellaCacheArbiter_covSum <= HellaCacheArbiter_covSum + 1'h1;
    end
  end
  always @(posedge clock) begin
    if(HellaCacheArbiter_cov_write_en & HellaCacheArbiter_cov_write_mask) begin
      HellaCacheArbiter_cov[HellaCacheArbiter_cov_write_addr] <= HellaCacheArbiter_cov_write_data; // @[Coverage map for HellaCacheArbiter]
    end
  end
endmodule
module PTW(
  input         clock,
  input         reset,
  output        io_requestor_0_req_ready,
  input         io_requestor_0_req_valid,
  input  [26:0] io_requestor_0_req_bits_bits_addr,
  output        io_requestor_0_resp_valid,
  output        io_requestor_0_resp_bits_ae,
  output [53:0] io_requestor_0_resp_bits_pte_ppn,
  output        io_requestor_0_resp_bits_pte_d,
  output        io_requestor_0_resp_bits_pte_a,
  output        io_requestor_0_resp_bits_pte_g,
  output        io_requestor_0_resp_bits_pte_u,
  output        io_requestor_0_resp_bits_pte_x,
  output        io_requestor_0_resp_bits_pte_w,
  output        io_requestor_0_resp_bits_pte_r,
  output        io_requestor_0_resp_bits_pte_v,
  output [1:0]  io_requestor_0_resp_bits_level,
  output        io_requestor_0_resp_bits_homogeneous,
  output [3:0]  io_requestor_0_ptbr_mode,
  output [1:0]  io_requestor_0_status_dprv,
  output        io_requestor_0_status_mxr,
  output        io_requestor_0_status_sum,
  output        io_requestor_0_pmp_0_cfg_l,
  output [1:0]  io_requestor_0_pmp_0_cfg_a,
  output        io_requestor_0_pmp_0_cfg_x,
  output        io_requestor_0_pmp_0_cfg_w,
  output        io_requestor_0_pmp_0_cfg_r,
  output [29:0] io_requestor_0_pmp_0_addr,
  output [31:0] io_requestor_0_pmp_0_mask,
  output        io_requestor_0_pmp_1_cfg_l,
  output [1:0]  io_requestor_0_pmp_1_cfg_a,
  output        io_requestor_0_pmp_1_cfg_x,
  output        io_requestor_0_pmp_1_cfg_w,
  output        io_requestor_0_pmp_1_cfg_r,
  output [29:0] io_requestor_0_pmp_1_addr,
  output [31:0] io_requestor_0_pmp_1_mask,
  output        io_requestor_0_pmp_2_cfg_l,
  output [1:0]  io_requestor_0_pmp_2_cfg_a,
  output        io_requestor_0_pmp_2_cfg_x,
  output        io_requestor_0_pmp_2_cfg_w,
  output        io_requestor_0_pmp_2_cfg_r,
  output [29:0] io_requestor_0_pmp_2_addr,
  output [31:0] io_requestor_0_pmp_2_mask,
  output        io_requestor_0_pmp_3_cfg_l,
  output [1:0]  io_requestor_0_pmp_3_cfg_a,
  output        io_requestor_0_pmp_3_cfg_x,
  output        io_requestor_0_pmp_3_cfg_w,
  output        io_requestor_0_pmp_3_cfg_r,
  output [29:0] io_requestor_0_pmp_3_addr,
  output [31:0] io_requestor_0_pmp_3_mask,
  output        io_requestor_0_pmp_4_cfg_l,
  output [1:0]  io_requestor_0_pmp_4_cfg_a,
  output        io_requestor_0_pmp_4_cfg_x,
  output        io_requestor_0_pmp_4_cfg_w,
  output        io_requestor_0_pmp_4_cfg_r,
  output [29:0] io_requestor_0_pmp_4_addr,
  output [31:0] io_requestor_0_pmp_4_mask,
  output        io_requestor_0_pmp_5_cfg_l,
  output [1:0]  io_requestor_0_pmp_5_cfg_a,
  output        io_requestor_0_pmp_5_cfg_x,
  output        io_requestor_0_pmp_5_cfg_w,
  output        io_requestor_0_pmp_5_cfg_r,
  output [29:0] io_requestor_0_pmp_5_addr,
  output [31:0] io_requestor_0_pmp_5_mask,
  output        io_requestor_0_pmp_6_cfg_l,
  output [1:0]  io_requestor_0_pmp_6_cfg_a,
  output        io_requestor_0_pmp_6_cfg_x,
  output        io_requestor_0_pmp_6_cfg_w,
  output        io_requestor_0_pmp_6_cfg_r,
  output [29:0] io_requestor_0_pmp_6_addr,
  output [31:0] io_requestor_0_pmp_6_mask,
  output        io_requestor_0_pmp_7_cfg_l,
  output [1:0]  io_requestor_0_pmp_7_cfg_a,
  output        io_requestor_0_pmp_7_cfg_x,
  output        io_requestor_0_pmp_7_cfg_w,
  output        io_requestor_0_pmp_7_cfg_r,
  output [29:0] io_requestor_0_pmp_7_addr,
  output [31:0] io_requestor_0_pmp_7_mask,
  output [26:0] io_requestor_0_vpoffset_bits_value,
  output        io_requestor_1_req_ready,
  input         io_requestor_1_req_valid,
  input         io_requestor_1_req_bits_valid,
  input  [26:0] io_requestor_1_req_bits_bits_addr,
  output        io_requestor_1_resp_valid,
  output        io_requestor_1_resp_bits_ae,
  output [53:0] io_requestor_1_resp_bits_pte_ppn,
  output        io_requestor_1_resp_bits_pte_d,
  output        io_requestor_1_resp_bits_pte_a,
  output        io_requestor_1_resp_bits_pte_g,
  output        io_requestor_1_resp_bits_pte_u,
  output        io_requestor_1_resp_bits_pte_x,
  output        io_requestor_1_resp_bits_pte_w,
  output        io_requestor_1_resp_bits_pte_r,
  output        io_requestor_1_resp_bits_pte_v,
  output [1:0]  io_requestor_1_resp_bits_level,
  output        io_requestor_1_resp_bits_homogeneous,
  output [3:0]  io_requestor_1_ptbr_mode,
  output [1:0]  io_requestor_1_status_prv,
  output        io_requestor_1_pmp_0_cfg_l,
  output [1:0]  io_requestor_1_pmp_0_cfg_a,
  output        io_requestor_1_pmp_0_cfg_x,
  output        io_requestor_1_pmp_0_cfg_w,
  output        io_requestor_1_pmp_0_cfg_r,
  output [29:0] io_requestor_1_pmp_0_addr,
  output [31:0] io_requestor_1_pmp_0_mask,
  output        io_requestor_1_pmp_1_cfg_l,
  output [1:0]  io_requestor_1_pmp_1_cfg_a,
  output        io_requestor_1_pmp_1_cfg_x,
  output        io_requestor_1_pmp_1_cfg_w,
  output        io_requestor_1_pmp_1_cfg_r,
  output [29:0] io_requestor_1_pmp_1_addr,
  output [31:0] io_requestor_1_pmp_1_mask,
  output        io_requestor_1_pmp_2_cfg_l,
  output [1:0]  io_requestor_1_pmp_2_cfg_a,
  output        io_requestor_1_pmp_2_cfg_x,
  output        io_requestor_1_pmp_2_cfg_w,
  output        io_requestor_1_pmp_2_cfg_r,
  output [29:0] io_requestor_1_pmp_2_addr,
  output [31:0] io_requestor_1_pmp_2_mask,
  output        io_requestor_1_pmp_3_cfg_l,
  output [1:0]  io_requestor_1_pmp_3_cfg_a,
  output        io_requestor_1_pmp_3_cfg_x,
  output        io_requestor_1_pmp_3_cfg_w,
  output        io_requestor_1_pmp_3_cfg_r,
  output [29:0] io_requestor_1_pmp_3_addr,
  output [31:0] io_requestor_1_pmp_3_mask,
  output        io_requestor_1_pmp_4_cfg_l,
  output [1:0]  io_requestor_1_pmp_4_cfg_a,
  output        io_requestor_1_pmp_4_cfg_x,
  output        io_requestor_1_pmp_4_cfg_w,
  output        io_requestor_1_pmp_4_cfg_r,
  output [29:0] io_requestor_1_pmp_4_addr,
  output [31:0] io_requestor_1_pmp_4_mask,
  output        io_requestor_1_pmp_5_cfg_l,
  output [1:0]  io_requestor_1_pmp_5_cfg_a,
  output        io_requestor_1_pmp_5_cfg_x,
  output        io_requestor_1_pmp_5_cfg_w,
  output        io_requestor_1_pmp_5_cfg_r,
  output [29:0] io_requestor_1_pmp_5_addr,
  output [31:0] io_requestor_1_pmp_5_mask,
  output        io_requestor_1_pmp_6_cfg_l,
  output [1:0]  io_requestor_1_pmp_6_cfg_a,
  output        io_requestor_1_pmp_6_cfg_x,
  output        io_requestor_1_pmp_6_cfg_w,
  output        io_requestor_1_pmp_6_cfg_r,
  output [29:0] io_requestor_1_pmp_6_addr,
  output [31:0] io_requestor_1_pmp_6_mask,
  output        io_requestor_1_pmp_7_cfg_l,
  output [1:0]  io_requestor_1_pmp_7_cfg_a,
  output        io_requestor_1_pmp_7_cfg_x,
  output        io_requestor_1_pmp_7_cfg_w,
  output        io_requestor_1_pmp_7_cfg_r,
  output [29:0] io_requestor_1_pmp_7_addr,
  output [31:0] io_requestor_1_pmp_7_mask,
  output [26:0] io_requestor_1_vpoffset_bits_value,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [39:0] io_mem_req_bits_addr,
  output        io_mem_s1_kill,
  input         io_mem_s2_nack,
  input         io_mem_resp_valid,
  input  [63:0] io_mem_resp_bits_data_word_bypass,
  input         io_mem_s2_xcpt_ae_ld,
  input  [3:0]  io_dpath_ptbr_mode,
  input  [43:0] io_dpath_ptbr_ppn,
  input         io_dpath_sfence_valid,
  input         io_dpath_sfence_bits_rs1,
  input  [1:0]  io_dpath_status_dprv,
  input  [1:0]  io_dpath_status_prv,
  input         io_dpath_status_mxr,
  input         io_dpath_status_sum,
  input         io_dpath_pmp_0_cfg_l,
  input  [1:0]  io_dpath_pmp_0_cfg_a,
  input         io_dpath_pmp_0_cfg_x,
  input         io_dpath_pmp_0_cfg_w,
  input         io_dpath_pmp_0_cfg_r,
  input  [29:0] io_dpath_pmp_0_addr,
  input  [31:0] io_dpath_pmp_0_mask,
  input         io_dpath_pmp_1_cfg_l,
  input  [1:0]  io_dpath_pmp_1_cfg_a,
  input         io_dpath_pmp_1_cfg_x,
  input         io_dpath_pmp_1_cfg_w,
  input         io_dpath_pmp_1_cfg_r,
  input  [29:0] io_dpath_pmp_1_addr,
  input  [31:0] io_dpath_pmp_1_mask,
  input         io_dpath_pmp_2_cfg_l,
  input  [1:0]  io_dpath_pmp_2_cfg_a,
  input         io_dpath_pmp_2_cfg_x,
  input         io_dpath_pmp_2_cfg_w,
  input         io_dpath_pmp_2_cfg_r,
  input  [29:0] io_dpath_pmp_2_addr,
  input  [31:0] io_dpath_pmp_2_mask,
  input         io_dpath_pmp_3_cfg_l,
  input  [1:0]  io_dpath_pmp_3_cfg_a,
  input         io_dpath_pmp_3_cfg_x,
  input         io_dpath_pmp_3_cfg_w,
  input         io_dpath_pmp_3_cfg_r,
  input  [29:0] io_dpath_pmp_3_addr,
  input  [31:0] io_dpath_pmp_3_mask,
  input         io_dpath_pmp_4_cfg_l,
  input  [1:0]  io_dpath_pmp_4_cfg_a,
  input         io_dpath_pmp_4_cfg_x,
  input         io_dpath_pmp_4_cfg_w,
  input         io_dpath_pmp_4_cfg_r,
  input  [29:0] io_dpath_pmp_4_addr,
  input  [31:0] io_dpath_pmp_4_mask,
  input         io_dpath_pmp_5_cfg_l,
  input  [1:0]  io_dpath_pmp_5_cfg_a,
  input         io_dpath_pmp_5_cfg_x,
  input         io_dpath_pmp_5_cfg_w,
  input         io_dpath_pmp_5_cfg_r,
  input  [29:0] io_dpath_pmp_5_addr,
  input  [31:0] io_dpath_pmp_5_mask,
  input         io_dpath_pmp_6_cfg_l,
  input  [1:0]  io_dpath_pmp_6_cfg_a,
  input         io_dpath_pmp_6_cfg_x,
  input         io_dpath_pmp_6_cfg_w,
  input         io_dpath_pmp_6_cfg_r,
  input  [29:0] io_dpath_pmp_6_addr,
  input  [31:0] io_dpath_pmp_6_mask,
  input         io_dpath_pmp_7_cfg_l,
  input  [1:0]  io_dpath_pmp_7_cfg_a,
  input         io_dpath_pmp_7_cfg_x,
  input         io_dpath_pmp_7_cfg_w,
  input         io_dpath_pmp_7_cfg_r,
  input  [29:0] io_dpath_pmp_7_addr,
  input  [31:0] io_dpath_pmp_7_mask,
  input         io_dpath_pcode_req_valid,
  input  [1:0]  io_dpath_pcode_req_bits_id,
  input  [19:0] io_dpath_pcode_req_bits_value_base,
  input  [9:0]  io_dpath_pcode_req_bits_value_mask,
  input         io_dpath_pcode_req_bits_value_valid,
  input         io_dpath_pcode_req_bits_value_locked,
  input  [26:0] io_dpath_vpoffset_req_bits_value,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         arb_halt
);
  wire  arb_clock; // @[PTW.scala 197:19]
  wire  arb_io_in_0_ready; // @[PTW.scala 197:19]
  wire  arb_io_in_0_valid; // @[PTW.scala 197:19]
  wire [26:0] arb_io_in_0_bits_bits_addr; // @[PTW.scala 197:19]
  wire  arb_io_in_1_ready; // @[PTW.scala 197:19]
  wire  arb_io_in_1_valid; // @[PTW.scala 197:19]
  wire  arb_io_in_1_bits_valid; // @[PTW.scala 197:19]
  wire [26:0] arb_io_in_1_bits_bits_addr; // @[PTW.scala 197:19]
  wire  arb_io_out_ready; // @[PTW.scala 197:19]
  wire  arb_io_out_valid; // @[PTW.scala 197:19]
  wire  arb_io_out_bits_valid; // @[PTW.scala 197:19]
  wire [26:0] arb_io_out_bits_bits_addr; // @[PTW.scala 197:19]
  wire  arb_io_chosen; // @[PTW.scala 197:19]
  wire [29:0] arb_io_covSum; // @[PTW.scala 197:19]
  wire  arb_metaAssert; // @[PTW.scala 197:19]
  wire  arb_metaReset; // @[PTW.scala 197:19]
  wire [53:0] pCodeLock_io_in_ppn; // @[PTW.scala 431:25]
  wire [1:0] pCodeLock_io_in_reserved_for_software; // @[PTW.scala 431:25]
  wire  pCodeLock_io_in_d; // @[PTW.scala 431:25]
  wire  pCodeLock_io_in_a; // @[PTW.scala 431:25]
  wire  pCodeLock_io_in_g; // @[PTW.scala 431:25]
  wire  pCodeLock_io_in_u; // @[PTW.scala 431:25]
  wire  pCodeLock_io_in_x; // @[PTW.scala 431:25]
  wire  pCodeLock_io_in_w; // @[PTW.scala 431:25]
  wire  pCodeLock_io_in_r; // @[PTW.scala 431:25]
  wire  pCodeLock_io_in_v; // @[PTW.scala 431:25]
  wire [53:0] pCodeLock_io_out_ppn; // @[PTW.scala 431:25]
  wire [1:0] pCodeLock_io_out_reserved_for_software; // @[PTW.scala 431:25]
  wire  pCodeLock_io_out_d; // @[PTW.scala 431:25]
  wire  pCodeLock_io_out_a; // @[PTW.scala 431:25]
  wire  pCodeLock_io_out_g; // @[PTW.scala 431:25]
  wire  pCodeLock_io_out_u; // @[PTW.scala 431:25]
  wire  pCodeLock_io_out_x; // @[PTW.scala 431:25]
  wire  pCodeLock_io_out_w; // @[PTW.scala 431:25]
  wire  pCodeLock_io_out_r; // @[PTW.scala 431:25]
  wire  pCodeLock_io_out_v; // @[PTW.scala 431:25]
  wire [19:0] pCodeLock_io_cfg_0_base; // @[PTW.scala 431:25]
  wire [9:0] pCodeLock_io_cfg_0_mask; // @[PTW.scala 431:25]
  wire  pCodeLock_io_cfg_0_valid; // @[PTW.scala 431:25]
  wire  pCodeLock_io_cfg_0_enable; // @[PTW.scala 431:25]
  wire [19:0] pCodeLock_io_cfg_1_base; // @[PTW.scala 431:25]
  wire [9:0] pCodeLock_io_cfg_1_mask; // @[PTW.scala 431:25]
  wire  pCodeLock_io_cfg_1_valid; // @[PTW.scala 431:25]
  wire  pCodeLock_io_cfg_1_enable; // @[PTW.scala 431:25]
  wire [19:0] pCodeLock_io_cfg_2_base; // @[PTW.scala 431:25]
  wire [9:0] pCodeLock_io_cfg_2_mask; // @[PTW.scala 431:25]
  wire  pCodeLock_io_cfg_2_valid; // @[PTW.scala 431:25]
  wire  pCodeLock_io_cfg_2_enable; // @[PTW.scala 431:25]
  wire [19:0] pCodeLock_io_cfg_3_base; // @[PTW.scala 431:25]
  wire [9:0] pCodeLock_io_cfg_3_mask; // @[PTW.scala 431:25]
  wire  pCodeLock_io_cfg_3_valid; // @[PTW.scala 431:25]
  wire  pCodeLock_io_cfg_3_enable; // @[PTW.scala 431:25]
  wire [29:0] pCodeLock_io_covSum; // @[PTW.scala 431:25]
  wire  pCodeLock_metaAssert; // @[PTW.scala 431:25]
  reg [19:0] pcode_cfg_0_base; // @[PTW.scala 160:22]
  reg [31:0] _RAND_0;
  reg [9:0] pcode_cfg_0_mask; // @[PTW.scala 160:22]
  reg [31:0] _RAND_1;
  reg  pcode_cfg_0_valid; // @[PTW.scala 160:22]
  reg [31:0] _RAND_2;
  reg  pcode_cfg_0_enable; // @[PTW.scala 160:22]
  reg [31:0] _RAND_3;
  reg [19:0] pcode_cfg_1_base; // @[PTW.scala 160:22]
  reg [31:0] _RAND_4;
  reg [9:0] pcode_cfg_1_mask; // @[PTW.scala 160:22]
  reg [31:0] _RAND_5;
  reg  pcode_cfg_1_valid; // @[PTW.scala 160:22]
  reg [31:0] _RAND_6;
  reg  pcode_cfg_1_enable; // @[PTW.scala 160:22]
  reg [31:0] _RAND_7;
  reg [19:0] pcode_cfg_2_base; // @[PTW.scala 160:22]
  reg [31:0] _RAND_8;
  reg [9:0] pcode_cfg_2_mask; // @[PTW.scala 160:22]
  reg [31:0] _RAND_9;
  reg  pcode_cfg_2_valid; // @[PTW.scala 160:22]
  reg [31:0] _RAND_10;
  reg  pcode_cfg_2_enable; // @[PTW.scala 160:22]
  reg [31:0] _RAND_11;
  reg [19:0] pcode_cfg_3_base; // @[PTW.scala 160:22]
  reg [31:0] _RAND_12;
  reg [9:0] pcode_cfg_3_mask; // @[PTW.scala 160:22]
  reg [31:0] _RAND_13;
  reg  pcode_cfg_3_valid; // @[PTW.scala 160:22]
  reg [31:0] _RAND_14;
  reg  pcode_cfg_3_enable; // @[PTW.scala 160:22]
  reg [31:0] _RAND_15;
  reg [2:0] state; // @[PTW.scala 195:18]
  reg [31:0] _RAND_16;
  reg  resp_valid_0; // @[PTW.scala 201:23]
  reg [31:0] _RAND_17;
  reg  resp_valid_1; // @[PTW.scala 201:23]
  reg [31:0] _RAND_18;
  wire  _T_582; // @[PTW.scala 202:24]
  reg  invalidated; // @[PTW.scala 208:24]
  reg [31:0] _RAND_19;
  reg [1:0] count; // @[PTW.scala 209:18]
  reg [31:0] _RAND_20;
  reg  resp_ae; // @[PTW.scala 210:24]
  reg [31:0] _RAND_21;
  reg [26:0] r_req_addr; // @[PTW.scala 213:18]
  reg [31:0] _RAND_22;
  reg  r_req_dest; // @[PTW.scala 214:23]
  reg [31:0] _RAND_23;
  reg [53:0] r_pte_ppn; // @[PTW.scala 215:18]
  reg [63:0] _RAND_24;
  reg [1:0] r_pte_reserved_for_software; // @[PTW.scala 215:18]
  reg [31:0] _RAND_25;
  reg  r_pte_d; // @[PTW.scala 215:18]
  reg [31:0] _RAND_26;
  reg  r_pte_a; // @[PTW.scala 215:18]
  reg [31:0] _RAND_27;
  reg  r_pte_g; // @[PTW.scala 215:18]
  reg [31:0] _RAND_28;
  reg  r_pte_u; // @[PTW.scala 215:18]
  reg [31:0] _RAND_29;
  reg  r_pte_x; // @[PTW.scala 215:18]
  reg [31:0] _RAND_30;
  reg  r_pte_w; // @[PTW.scala 215:18]
  reg [31:0] _RAND_31;
  reg  r_pte_r; // @[PTW.scala 215:18]
  reg [31:0] _RAND_32;
  reg  r_pte_v; // @[PTW.scala 215:18]
  reg [31:0] _RAND_33;
  wire  tmp_v; // @[PTW.scala 218:33]
  wire  tmp_r; // @[PTW.scala 218:33]
  wire  tmp_w; // @[PTW.scala 218:33]
  wire  tmp_x; // @[PTW.scala 218:33]
  wire  tmp_u; // @[PTW.scala 218:33]
  wire  tmp_g; // @[PTW.scala 218:33]
  wire  tmp_a; // @[PTW.scala 218:33]
  wire  tmp_d; // @[PTW.scala 218:33]
  wire [1:0] tmp_reserved_for_software; // @[PTW.scala 218:33]
  wire [53:0] tmp_ppn; // @[PTW.scala 218:33]
  wire  _T_624; // @[PTW.scala 221:17]
  wire  _T_625; // @[PTW.scala 221:26]
  wire  _T_626; // @[PTW.scala 224:21]
  wire  _T_628; // @[PTW.scala 224:95]
  wire  _T_629; // @[PTW.scala 224:26]
  wire  _GEN_37; // @[PTW.scala 224:102]
  wire  _T_630; // @[PTW.scala 224:21]
  wire  _T_632; // @[PTW.scala 224:95]
  wire  _T_633; // @[PTW.scala 224:26]
  wire  _GEN_38; // @[PTW.scala 224:102]
  wire  res_v; // @[PTW.scala 221:36]
  wire  invalid_paddr; // @[PTW.scala 226:32]
  wire  _T_636; // @[PTW.scala 76:33]
  wire  _T_638; // @[PTW.scala 76:39]
  wire  _T_640; // @[PTW.scala 76:45]
  wire  _T_642; // @[PTW.scala 228:30]
  wire  _T_643; // @[PTW.scala 228:57]
  wire  traverse; // @[PTW.scala 228:48]
  wire  _T_650; // @[package.scala 31:81]
  wire [8:0] _T_651; // @[package.scala 31:71]
  wire  _T_652; // @[package.scala 31:81]
  wire [8:0] _T_653; // @[package.scala 31:71]
  wire  _T_654; // @[package.scala 31:81]
  wire [8:0] vpn_idx; // @[package.scala 31:71]
  wire [62:0] _T_655; // @[Cat.scala 30:58]
  wire [65:0] pte_addr; // @[PTW.scala 232:29]
  wire [53:0] _T_658; // @[Cat.scala 30:58]
  wire [53:0] _T_661; // @[Cat.scala 30:58]
  wire [53:0] fragmented_superpage_ppn; // @[package.scala 31:71]
  wire  _T_665; // @[Decoupled.scala 37:37]
  reg [6:0] _T_667; // @[Replacement.scala 41:30]
  reg [31:0] _RAND_34;
  reg  invalid; // @[PTW.scala 247:26]
  reg [31:0] _RAND_35;
  reg [7:0] reg_valid; // @[PTW.scala 248:24]
  reg [31:0] _RAND_36;
  wire [7:0] valid; // @[PTW.scala 249:20]
  reg [31:0] tags_0; // @[PTW.scala 250:19]
  reg [31:0] _RAND_37;
  reg [31:0] tags_1; // @[PTW.scala 250:19]
  reg [31:0] _RAND_38;
  reg [31:0] tags_2; // @[PTW.scala 250:19]
  reg [31:0] _RAND_39;
  reg [31:0] tags_3; // @[PTW.scala 250:19]
  reg [31:0] _RAND_40;
  reg [31:0] tags_4; // @[PTW.scala 250:19]
  reg [31:0] _RAND_41;
  reg [31:0] tags_5; // @[PTW.scala 250:19]
  reg [31:0] _RAND_42;
  reg [31:0] tags_6; // @[PTW.scala 250:19]
  reg [31:0] _RAND_43;
  reg [31:0] tags_7; // @[PTW.scala 250:19]
  reg [31:0] _RAND_44;
  reg [19:0] data_0; // @[PTW.scala 251:19]
  reg [31:0] _RAND_45;
  reg [19:0] data_1; // @[PTW.scala 251:19]
  reg [31:0] _RAND_46;
  reg [19:0] data_2; // @[PTW.scala 251:19]
  reg [31:0] _RAND_47;
  reg [19:0] data_3; // @[PTW.scala 251:19]
  reg [31:0] _RAND_48;
  reg [19:0] data_4; // @[PTW.scala 251:19]
  reg [31:0] _RAND_49;
  reg [19:0] data_5; // @[PTW.scala 251:19]
  reg [31:0] _RAND_50;
  reg [19:0] data_6; // @[PTW.scala 251:19]
  reg [31:0] _RAND_51;
  reg [19:0] data_7; // @[PTW.scala 251:19]
  reg [31:0] _RAND_52;
  wire [65:0] _GEN_148; // @[PTW.scala 253:27]
  wire  _T_696; // @[PTW.scala 253:27]
  wire [65:0] _GEN_149; // @[PTW.scala 253:27]
  wire  _T_697; // @[PTW.scala 253:27]
  wire [65:0] _GEN_150; // @[PTW.scala 253:27]
  wire  _T_698; // @[PTW.scala 253:27]
  wire [65:0] _GEN_151; // @[PTW.scala 253:27]
  wire  _T_699; // @[PTW.scala 253:27]
  wire [65:0] _GEN_152; // @[PTW.scala 253:27]
  wire  _T_700; // @[PTW.scala 253:27]
  wire [65:0] _GEN_153; // @[PTW.scala 253:27]
  wire  _T_701; // @[PTW.scala 253:27]
  wire [65:0] _GEN_154; // @[PTW.scala 253:27]
  wire  _T_702; // @[PTW.scala 253:27]
  wire [65:0] _GEN_155; // @[PTW.scala 253:27]
  wire  _T_703; // @[PTW.scala 253:27]
  wire [7:0] _T_710; // @[Cat.scala 30:58]
  wire [7:0] hits; // @[PTW.scala 253:48]
  wire  hit; // @[PTW.scala 254:20]
  wire  _T_711; // @[PTW.scala 255:18]
  wire  _T_712; // @[PTW.scala 255:39]
  wire  _T_713; // @[PTW.scala 255:30]
  wire  _T_714; // @[PTW.scala 255:52]
  wire  _T_716; // @[PTW.scala 255:64]
  wire  _T_718; // @[PTW.scala 255:72]
  wire  _T_720; // @[PTW.scala 256:25]
  wire [7:0] _T_721; // @[Replacement.scala 57:31]
  wire [7:0] _T_725; // @[Replacement.scala 61:48]
  wire [1:0] _T_728; // @[Cat.scala 30:58]
  wire [7:0] _T_732; // @[Replacement.scala 61:48]
  wire [2:0] _T_735; // @[Cat.scala 30:58]
  wire [7:0] _T_739; // @[Replacement.scala 61:48]
  wire [3:0] _T_742; // @[Cat.scala 30:58]
  wire  _T_745; // @[OneHot.scala 39:40]
  wire  _T_746; // @[OneHot.scala 39:40]
  wire  _T_747; // @[OneHot.scala 39:40]
  wire  _T_748; // @[OneHot.scala 39:40]
  wire  _T_749; // @[OneHot.scala 39:40]
  wire  _T_750; // @[OneHot.scala 39:40]
  wire  _T_751; // @[OneHot.scala 39:40]
  wire [2:0] _T_753; // @[Mux.scala 31:69]
  wire [2:0] _T_754; // @[Mux.scala 31:69]
  wire [2:0] _T_755; // @[Mux.scala 31:69]
  wire [2:0] _T_756; // @[Mux.scala 31:69]
  wire [2:0] _T_757; // @[Mux.scala 31:69]
  wire [2:0] _T_758; // @[Mux.scala 31:69]
  wire [2:0] _T_759; // @[Mux.scala 31:69]
  wire [2:0] r; // @[PTW.scala 256:18]
  wire [7:0] _T_760; // @[OneHot.scala 45:35]
  wire [7:0] _T_761; // @[PTW.scala 258:49]
  wire [7:0] _T_764; // @[PTW.scala 258:70]
  wire [53:0] res_ppn; // @[PTW.scala 220:13]
  wire  _GEN_58; // @[PTW.scala 255:89]
  wire  _T_768; // @[PTW.scala 262:24]
  wire  _T_769; // @[PTW.scala 262:15]
  wire  _T_772; // @[OneHot.scala 28:14]
  wire [3:0] _T_773; // @[OneHot.scala 28:28]
  wire  _T_776; // @[OneHot.scala 28:14]
  wire [1:0] _T_777; // @[OneHot.scala 28:28]
  wire [2:0] _T_780; // @[Cat.scala 30:58]
  wire [7:0] _T_785; // @[Replacement.scala 50:37]
  wire [7:0] _T_787; // @[Replacement.scala 50:37]
  wire [7:0] _T_789; // @[Replacement.scala 50:37]
  wire [1:0] _T_790; // @[Cat.scala 30:58]
  wire [3:0] _T_793; // @[Replacement.scala 50:37]
  wire [7:0] _GEN_157; // @[Replacement.scala 50:37]
  wire [7:0] _T_794; // @[Replacement.scala 50:37]
  wire [7:0] _T_796; // @[Replacement.scala 50:37]
  wire [7:0] _T_798; // @[Replacement.scala 50:37]
  wire [2:0] _T_799; // @[Cat.scala 30:58]
  wire [7:0] _T_802; // @[Replacement.scala 50:37]
  wire [7:0] _T_803; // @[Replacement.scala 50:37]
  wire [7:0] _T_805; // @[Replacement.scala 50:37]
  wire [7:0] _T_807; // @[Replacement.scala 50:37]
  wire  _T_811; // @[PTW.scala 263:33]
  wire  _GEN_77; // @[PTW.scala 263:63]
  wire  pte_cache_hit; // @[PTW.scala 268:10]
  wire [19:0] _T_830; // @[Mux.scala 19:72]
  wire [19:0] _T_831; // @[Mux.scala 19:72]
  wire [19:0] _T_832; // @[Mux.scala 19:72]
  wire [19:0] _T_833; // @[Mux.scala 19:72]
  wire [19:0] _T_834; // @[Mux.scala 19:72]
  wire [19:0] _T_835; // @[Mux.scala 19:72]
  wire [19:0] _T_836; // @[Mux.scala 19:72]
  wire [19:0] _T_837; // @[Mux.scala 19:72]
  wire [19:0] _T_838; // @[Mux.scala 19:72]
  wire [19:0] _T_839; // @[Mux.scala 19:72]
  wire [19:0] _T_840; // @[Mux.scala 19:72]
  wire [19:0] _T_841; // @[Mux.scala 19:72]
  wire [19:0] _T_842; // @[Mux.scala 19:72]
  wire [19:0] _T_843; // @[Mux.scala 19:72]
  wire [19:0] pte_cache_data; // @[Mux.scala 19:72]
  wire  _T_849; // @[PTW.scala 341:56]
  wire  _T_852; // @[PTW.scala 343:48]
  wire [65:0] _T_862; // @[Parameters.scala 121:31]
  wire [66:0] _T_863; // @[Parameters.scala 121:49]
  wire [66:0] _T_865; // @[Parameters.scala 121:52]
  wire  _T_866; // @[Parameters.scala 121:67]
  wire [65:0] _T_867; // @[Parameters.scala 121:31]
  wire [66:0] _T_868; // @[Parameters.scala 121:49]
  wire [66:0] _T_870; // @[Parameters.scala 121:52]
  wire  _T_871; // @[Parameters.scala 121:67]
  wire [65:0] _T_872; // @[Parameters.scala 121:31]
  wire [66:0] _T_873; // @[Parameters.scala 121:49]
  wire [66:0] _T_875; // @[Parameters.scala 121:52]
  wire  _T_876; // @[Parameters.scala 121:67]
  wire  _T_878; // @[TLBPermissions.scala 97:65]
  wire  _T_879; // @[TLBPermissions.scala 97:65]
  wire [66:0] _T_883; // @[Parameters.scala 121:49]
  wire [65:0] _T_912; // @[Parameters.scala 121:31]
  wire [66:0] _T_913; // @[Parameters.scala 121:49]
  wire [66:0] _T_915; // @[Parameters.scala 121:52]
  wire  _T_916; // @[Parameters.scala 121:67]
  wire [65:0] _T_922; // @[Parameters.scala 121:31]
  wire [66:0] _T_923; // @[Parameters.scala 121:49]
  wire [66:0] _T_925; // @[Parameters.scala 121:52]
  wire  _T_926; // @[Parameters.scala 121:67]
  wire [65:0] _T_927; // @[Parameters.scala 121:31]
  wire [66:0] _T_928; // @[Parameters.scala 121:49]
  wire [66:0] _T_930; // @[Parameters.scala 121:52]
  wire  _T_931; // @[Parameters.scala 121:67]
  wire [66:0] _T_940; // @[Parameters.scala 121:52]
  wire  _T_941; // @[Parameters.scala 121:67]
  wire  _T_943; // @[TLBPermissions.scala 97:65]
  wire  _T_944; // @[TLBPermissions.scala 97:65]
  wire  _T_945; // @[TLBPermissions.scala 97:65]
  wire  _T_946; // @[TLBPermissions.scala 97:65]
  wire  _T_947; // @[TLBPermissions.scala 97:65]
  wire  _T_948; // @[TLBPermissions.scala 97:65]
  wire  _T_1001; // @[package.scala 31:71]
  wire  _T_1003; // @[package.scala 31:71]
  wire  pmaHomogeneous; // @[package.scala 31:71]
  wire [65:0] _T_1006; // @[PTW.scala 362:92]
  wire  _T_1025; // @[package.scala 31:71]
  wire  _T_1027; // @[package.scala 31:71]
  wire  _T_1029; // @[package.scala 31:71]
  wire [31:0] _T_1030; // @[PMP.scala 54:36]
  wire [31:0] _T_1032; // @[PMP.scala 54:48]
  wire [65:0] _GEN_159; // @[PMP.scala 92:53]
  wire [65:0] _T_1034; // @[PMP.scala 92:53]
  wire  _T_1036; // @[PMP.scala 92:78]
  wire  _T_1043; // @[PMP.scala 92:78]
  wire  _T_1050; // @[PMP.scala 92:78]
  wire  _T_1052; // @[package.scala 31:71]
  wire  _T_1054; // @[package.scala 31:71]
  wire  _T_1056; // @[package.scala 31:71]
  wire  _T_1057; // @[PMP.scala 92:21]
  wire  _T_1070; // @[PMP.scala 101:32]
  wire [31:0] _T_1073; // @[package.scala 31:71]
  wire [31:0] _T_1075; // @[package.scala 31:71]
  wire [31:0] _T_1077; // @[package.scala 31:71]
  wire [65:0] _GEN_163; // @[PMP.scala 104:30]
  wire [65:0] _T_1078; // @[PMP.scala 104:30]
  wire [31:0] _T_1090; // @[PMP.scala 105:53]
  wire [65:0] _GEN_165; // @[PMP.scala 105:40]
  wire  _T_1091; // @[PMP.scala 105:40]
  wire  _T_1094; // @[PMP.scala 107:41]
  wire  _T_1095; // @[PMP.scala 112:58]
  wire  _T_1096; // @[PMP.scala 112:8]
  wire  _T_1103; // @[package.scala 31:71]
  wire  _T_1105; // @[package.scala 31:71]
  wire  _T_1107; // @[package.scala 31:71]
  wire [31:0] _T_1108; // @[PMP.scala 54:36]
  wire [31:0] _T_1110; // @[PMP.scala 54:48]
  wire [65:0] _GEN_166; // @[PMP.scala 92:53]
  wire [65:0] _T_1112; // @[PMP.scala 92:53]
  wire  _T_1114; // @[PMP.scala 92:78]
  wire  _T_1121; // @[PMP.scala 92:78]
  wire  _T_1128; // @[PMP.scala 92:78]
  wire  _T_1130; // @[package.scala 31:71]
  wire  _T_1132; // @[package.scala 31:71]
  wire  _T_1134; // @[package.scala 31:71]
  wire  _T_1135; // @[PMP.scala 92:21]
  wire  _T_1148; // @[PMP.scala 101:32]
  wire [31:0] _T_1168; // @[PMP.scala 105:53]
  wire [65:0] _GEN_174; // @[PMP.scala 105:40]
  wire  _T_1169; // @[PMP.scala 105:40]
  wire  _T_1170; // @[PMP.scala 107:21]
  wire  _T_1171; // @[PMP.scala 107:62]
  wire  _T_1172; // @[PMP.scala 107:41]
  wire  _T_1173; // @[PMP.scala 112:58]
  wire  _T_1174; // @[PMP.scala 112:8]
  wire  _T_1175; // @[PMP.scala 132:10]
  wire  _T_1181; // @[package.scala 31:71]
  wire  _T_1183; // @[package.scala 31:71]
  wire  _T_1185; // @[package.scala 31:71]
  wire [31:0] _T_1186; // @[PMP.scala 54:36]
  wire [31:0] _T_1188; // @[PMP.scala 54:48]
  wire [65:0] _GEN_175; // @[PMP.scala 92:53]
  wire [65:0] _T_1190; // @[PMP.scala 92:53]
  wire  _T_1192; // @[PMP.scala 92:78]
  wire  _T_1199; // @[PMP.scala 92:78]
  wire  _T_1206; // @[PMP.scala 92:78]
  wire  _T_1208; // @[package.scala 31:71]
  wire  _T_1210; // @[package.scala 31:71]
  wire  _T_1212; // @[package.scala 31:71]
  wire  _T_1213; // @[PMP.scala 92:21]
  wire  _T_1226; // @[PMP.scala 101:32]
  wire [31:0] _T_1246; // @[PMP.scala 105:53]
  wire [65:0] _GEN_183; // @[PMP.scala 105:40]
  wire  _T_1247; // @[PMP.scala 105:40]
  wire  _T_1248; // @[PMP.scala 107:21]
  wire  _T_1249; // @[PMP.scala 107:62]
  wire  _T_1250; // @[PMP.scala 107:41]
  wire  _T_1251; // @[PMP.scala 112:58]
  wire  _T_1252; // @[PMP.scala 112:8]
  wire  _T_1253; // @[PMP.scala 132:10]
  wire  _T_1259; // @[package.scala 31:71]
  wire  _T_1261; // @[package.scala 31:71]
  wire  _T_1263; // @[package.scala 31:71]
  wire [31:0] _T_1264; // @[PMP.scala 54:36]
  wire [31:0] _T_1266; // @[PMP.scala 54:48]
  wire [65:0] _GEN_184; // @[PMP.scala 92:53]
  wire [65:0] _T_1268; // @[PMP.scala 92:53]
  wire  _T_1270; // @[PMP.scala 92:78]
  wire  _T_1277; // @[PMP.scala 92:78]
  wire  _T_1284; // @[PMP.scala 92:78]
  wire  _T_1286; // @[package.scala 31:71]
  wire  _T_1288; // @[package.scala 31:71]
  wire  _T_1290; // @[package.scala 31:71]
  wire  _T_1291; // @[PMP.scala 92:21]
  wire  _T_1304; // @[PMP.scala 101:32]
  wire [31:0] _T_1324; // @[PMP.scala 105:53]
  wire [65:0] _GEN_192; // @[PMP.scala 105:40]
  wire  _T_1325; // @[PMP.scala 105:40]
  wire  _T_1326; // @[PMP.scala 107:21]
  wire  _T_1327; // @[PMP.scala 107:62]
  wire  _T_1328; // @[PMP.scala 107:41]
  wire  _T_1329; // @[PMP.scala 112:58]
  wire  _T_1330; // @[PMP.scala 112:8]
  wire  _T_1331; // @[PMP.scala 132:10]
  wire  _T_1337; // @[package.scala 31:71]
  wire  _T_1339; // @[package.scala 31:71]
  wire  _T_1341; // @[package.scala 31:71]
  wire [31:0] _T_1342; // @[PMP.scala 54:36]
  wire [31:0] _T_1344; // @[PMP.scala 54:48]
  wire [65:0] _GEN_193; // @[PMP.scala 92:53]
  wire [65:0] _T_1346; // @[PMP.scala 92:53]
  wire  _T_1348; // @[PMP.scala 92:78]
  wire  _T_1355; // @[PMP.scala 92:78]
  wire  _T_1362; // @[PMP.scala 92:78]
  wire  _T_1364; // @[package.scala 31:71]
  wire  _T_1366; // @[package.scala 31:71]
  wire  _T_1368; // @[package.scala 31:71]
  wire  _T_1369; // @[PMP.scala 92:21]
  wire  _T_1382; // @[PMP.scala 101:32]
  wire [31:0] _T_1402; // @[PMP.scala 105:53]
  wire [65:0] _GEN_201; // @[PMP.scala 105:40]
  wire  _T_1403; // @[PMP.scala 105:40]
  wire  _T_1404; // @[PMP.scala 107:21]
  wire  _T_1405; // @[PMP.scala 107:62]
  wire  _T_1406; // @[PMP.scala 107:41]
  wire  _T_1407; // @[PMP.scala 112:58]
  wire  _T_1408; // @[PMP.scala 112:8]
  wire  _T_1409; // @[PMP.scala 132:10]
  wire  _T_1415; // @[package.scala 31:71]
  wire  _T_1417; // @[package.scala 31:71]
  wire  _T_1419; // @[package.scala 31:71]
  wire [31:0] _T_1420; // @[PMP.scala 54:36]
  wire [31:0] _T_1422; // @[PMP.scala 54:48]
  wire [65:0] _GEN_202; // @[PMP.scala 92:53]
  wire [65:0] _T_1424; // @[PMP.scala 92:53]
  wire  _T_1426; // @[PMP.scala 92:78]
  wire  _T_1433; // @[PMP.scala 92:78]
  wire  _T_1440; // @[PMP.scala 92:78]
  wire  _T_1442; // @[package.scala 31:71]
  wire  _T_1444; // @[package.scala 31:71]
  wire  _T_1446; // @[package.scala 31:71]
  wire  _T_1447; // @[PMP.scala 92:21]
  wire  _T_1460; // @[PMP.scala 101:32]
  wire [31:0] _T_1480; // @[PMP.scala 105:53]
  wire [65:0] _GEN_210; // @[PMP.scala 105:40]
  wire  _T_1481; // @[PMP.scala 105:40]
  wire  _T_1482; // @[PMP.scala 107:21]
  wire  _T_1483; // @[PMP.scala 107:62]
  wire  _T_1484; // @[PMP.scala 107:41]
  wire  _T_1485; // @[PMP.scala 112:58]
  wire  _T_1486; // @[PMP.scala 112:8]
  wire  _T_1487; // @[PMP.scala 132:10]
  wire  _T_1493; // @[package.scala 31:71]
  wire  _T_1495; // @[package.scala 31:71]
  wire  _T_1497; // @[package.scala 31:71]
  wire [31:0] _T_1498; // @[PMP.scala 54:36]
  wire [31:0] _T_1500; // @[PMP.scala 54:48]
  wire [65:0] _GEN_211; // @[PMP.scala 92:53]
  wire [65:0] _T_1502; // @[PMP.scala 92:53]
  wire  _T_1504; // @[PMP.scala 92:78]
  wire  _T_1511; // @[PMP.scala 92:78]
  wire  _T_1518; // @[PMP.scala 92:78]
  wire  _T_1520; // @[package.scala 31:71]
  wire  _T_1522; // @[package.scala 31:71]
  wire  _T_1524; // @[package.scala 31:71]
  wire  _T_1525; // @[PMP.scala 92:21]
  wire  _T_1538; // @[PMP.scala 101:32]
  wire [31:0] _T_1558; // @[PMP.scala 105:53]
  wire [65:0] _GEN_219; // @[PMP.scala 105:40]
  wire  _T_1559; // @[PMP.scala 105:40]
  wire  _T_1560; // @[PMP.scala 107:21]
  wire  _T_1561; // @[PMP.scala 107:62]
  wire  _T_1562; // @[PMP.scala 107:41]
  wire  _T_1563; // @[PMP.scala 112:58]
  wire  _T_1564; // @[PMP.scala 112:8]
  wire  _T_1565; // @[PMP.scala 132:10]
  wire  _T_1571; // @[package.scala 31:71]
  wire  _T_1573; // @[package.scala 31:71]
  wire  _T_1575; // @[package.scala 31:71]
  wire [31:0] _T_1576; // @[PMP.scala 54:36]
  wire [31:0] _T_1578; // @[PMP.scala 54:48]
  wire [65:0] _GEN_220; // @[PMP.scala 92:53]
  wire [65:0] _T_1580; // @[PMP.scala 92:53]
  wire  _T_1582; // @[PMP.scala 92:78]
  wire  _T_1589; // @[PMP.scala 92:78]
  wire  _T_1596; // @[PMP.scala 92:78]
  wire  _T_1598; // @[package.scala 31:71]
  wire  _T_1600; // @[package.scala 31:71]
  wire  _T_1602; // @[package.scala 31:71]
  wire  _T_1603; // @[PMP.scala 92:21]
  wire  _T_1616; // @[PMP.scala 101:32]
  wire [31:0] _T_1636; // @[PMP.scala 105:53]
  wire [65:0] _GEN_228; // @[PMP.scala 105:40]
  wire  _T_1637; // @[PMP.scala 105:40]
  wire  _T_1638; // @[PMP.scala 107:21]
  wire  _T_1639; // @[PMP.scala 107:62]
  wire  _T_1640; // @[PMP.scala 107:41]
  wire  _T_1641; // @[PMP.scala 112:58]
  wire  _T_1642; // @[PMP.scala 112:8]
  wire  pmpHomogeneous; // @[PMP.scala 132:10]
  wire  homogeneous; // @[PTW.scala 363:36]
  wire  ae; // @[PTW.scala 492:22]
  wire [2:0] _GEN_136; // @[PTW.scala 487:21]
  wire  _T_1650; // @[Conditional.scala 37:30]
  wire [2:0] _T_1652; // @[PTW.scala 393:26]
  wire [2:0] _GEN_80; // @[PTW.scala 392:32]
  wire  _T_1653; // @[Conditional.scala 37:30]
  wire [2:0] _T_1656; // @[PTW.scala 401:26]
  wire [2:0] _GEN_82; // @[PTW.scala 398:28]
  wire  _T_1657; // @[Conditional.scala 37:30]
  wire  _T_1658; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_86; // @[PTW.scala 409:35]
  wire  _T_1664; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_93; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_99; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_105; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_112; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_117; // @[Conditional.scala 40:58]
  wire [2:0] _GEN_130; // @[PTW.scala 481:25]
  wire [2:0] next_state; // @[PTW.scala 485:28]
  wire [1:0] _T_1655; // @[PTW.scala 399:24]
  wire  _GEN_87; // @[PTW.scala 409:35]
  wire  _GEN_88; // @[PTW.scala 409:35]
  wire  _GEN_94; // @[Conditional.scala 39:67]
  wire  _GEN_95; // @[Conditional.scala 39:67]
  wire  _GEN_100; // @[Conditional.scala 39:67]
  wire  _GEN_101; // @[Conditional.scala 39:67]
  wire  _GEN_102; // @[Conditional.scala 39:67]
  wire  _GEN_107; // @[Conditional.scala 39:67]
  wire  _GEN_108; // @[Conditional.scala 39:67]
  wire  _GEN_114; // @[Conditional.scala 39:67]
  wire  _GEN_115; // @[Conditional.scala 39:67]
  wire  _GEN_120; // @[Conditional.scala 40:58]
  wire  _GEN_121; // @[Conditional.scala 40:58]
  wire  _T_1671; // @[PTW.scala 465:15]
  wire  _T_1673; // @[PTW.scala 465:40]
  wire  _T_1676; // @[PTW.scala 466:25]
  wire [53:0] pte_2_ppn; // @[PTW.scala 428:13]
  wire [53:0] _T_1680_ppn; // @[PTW.scala 467:8]
  wire [53:0] pte_1_ppn; // @[PTW.scala 428:13]
  wire [53:0] _T_1681_ppn; // @[PTW.scala 466:8]
  wire [1:0] _T_1681_reserved_for_software; // @[PTW.scala 466:8]
  wire  _T_1681_d; // @[PTW.scala 466:8]
  wire  _T_1681_a; // @[PTW.scala 466:8]
  wire  _T_1681_g; // @[PTW.scala 466:8]
  wire  _T_1681_u; // @[PTW.scala 466:8]
  wire  _T_1681_x; // @[PTW.scala 466:8]
  wire  _T_1681_w; // @[PTW.scala 466:8]
  wire  _T_1681_r; // @[PTW.scala 466:8]
  wire  _T_1681_v; // @[PTW.scala 466:8]
  wire [53:0] _T_1682_ppn; // @[PTW.scala 465:8]
  wire [1:0] _T_1682_reserved_for_software; // @[PTW.scala 465:8]
  wire  _T_1682_d; // @[PTW.scala 465:8]
  wire  _T_1682_a; // @[PTW.scala 465:8]
  wire  _T_1682_g; // @[PTW.scala 465:8]
  wire  _T_1682_u; // @[PTW.scala 465:8]
  wire  _T_1682_x; // @[PTW.scala 465:8]
  wire  _T_1682_w; // @[PTW.scala 465:8]
  wire  _T_1682_r; // @[PTW.scala 465:8]
  wire  _T_1682_v; // @[PTW.scala 465:8]
  wire [53:0] _T_1684_ppn; // @[PTW.scala 463:8]
  wire [1:0] _T_1684_reserved_for_software; // @[PTW.scala 463:8]
  wire  _T_1684_d; // @[PTW.scala 463:8]
  wire  _T_1684_a; // @[PTW.scala 463:8]
  wire  _T_1684_g; // @[PTW.scala 463:8]
  wire  _T_1684_u; // @[PTW.scala 463:8]
  wire  _T_1684_x; // @[PTW.scala 463:8]
  wire  _T_1684_w; // @[PTW.scala 463:8]
  wire  _T_1684_r; // @[PTW.scala 463:8]
  wire  _T_1684_v; // @[PTW.scala 463:8]
  wire [63:0] _T_1693; // @[package.scala 208:71]
  wire  _GEN_123; // @[PTW.scala 477:28]
  wire  _GEN_124; // @[PTW.scala 477:28]
  wire  _T_1723; // @[PTW.scala 482:11]
  wire  _T_1729; // @[PTW.scala 486:11]
  reg [19:0] PTW_state; // @[Register tracking PTW state]
  reg [31:0] _RAND_53;
  reg  PTW_cov [0:1048575]; // @[Coverage map for PTW]
  reg [31:0] _RAND_54;
  wire  PTW_cov_read_data; // @[Coverage map for PTW]
  wire [19:0] PTW_cov_read_addr; // @[Coverage map for PTW]
  wire  PTW_cov_write_data; // @[Coverage map for PTW]
  wire [19:0] PTW_cov_write_addr; // @[Coverage map for PTW]
  wire  PTW_cov_write_mask; // @[Coverage map for PTW]
  wire  PTW_cov_write_en; // @[Coverage map for PTW]
  reg [29:0] PTW_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_55;
  wire [16:0] count_shl;
  wire [19:0] count_pad;
  wire [10:0] invalid_shl;
  wire [19:0] invalid_pad;
  wire [10:0] state_shl;
  wire [19:0] state_pad;
  wire [9:0] reg_valid_shl;
  wire [19:0] reg_valid_pad;
  wire [9:0] _T_667_shl;
  wire [19:0] _T_667_pad;
  wire [8:0] invalidated_shl;
  wire [19:0] invalidated_pad;
  wire [12:0] pcode_cfg_0_enable_shl;
  wire [19:0] pcode_cfg_0_enable_pad;
  wire [19:0] pcode_cfg_0_base_shl;
  wire [19:0] pcode_cfg_0_base_pad;
  wire [15:0] pcode_cfg_0_mask_shl;
  wire [19:0] pcode_cfg_0_mask_pad;
  wire [1:0] pcode_cfg_0_valid_shl;
  wire [19:0] pcode_cfg_0_valid_pad;
  wire [19:0] PTW_xor3;
  wire [19:0] PTW_xor10;
  wire [19:0] PTW_xor4;
  wire [19:0] PTW_xor1;
  wire [19:0] PTW_xor5;
  wire [19:0] PTW_xor14;
  wire [19:0] PTW_xor6;
  wire [19:0] PTW_xor2;
  wire [19:0] PTW_xor0;
  wire [29:0] arb_sum;
  wire [29:0] pCodeLock_sum;
  wire  stopEn0;
  wire  stopEn1;
  wire  arb_metaAssert_wire;
  wire  pCodeLock_metaAssert_wire;
  wire  PTW_or1;
  wire  PTW_or2;
  wire  PTW_or0;
  reg  PTW_metaAssert;
  reg [31:0] _RAND_56;
  RRArbiter arb ( // @[PTW.scala 197:19]
    .clock(arb_clock),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_bits_addr(arb_io_in_0_bits_bits_addr),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_valid(arb_io_in_1_bits_valid),
    .io_in_1_bits_bits_addr(arb_io_in_1_bits_bits_addr),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_valid(arb_io_out_bits_valid),
    .io_out_bits_bits_addr(arb_io_out_bits_bits_addr),
    .io_chosen(arb_io_chosen),
    .io_covSum(arb_io_covSum),
    .metaAssert(arb_metaAssert),
    .metaReset(arb_metaReset)
  );
  PCodeLock pCodeLock ( // @[PTW.scala 431:25]
    .io_in_ppn(pCodeLock_io_in_ppn),
    .io_in_reserved_for_software(pCodeLock_io_in_reserved_for_software),
    .io_in_d(pCodeLock_io_in_d),
    .io_in_a(pCodeLock_io_in_a),
    .io_in_g(pCodeLock_io_in_g),
    .io_in_u(pCodeLock_io_in_u),
    .io_in_x(pCodeLock_io_in_x),
    .io_in_w(pCodeLock_io_in_w),
    .io_in_r(pCodeLock_io_in_r),
    .io_in_v(pCodeLock_io_in_v),
    .io_out_ppn(pCodeLock_io_out_ppn),
    .io_out_reserved_for_software(pCodeLock_io_out_reserved_for_software),
    .io_out_d(pCodeLock_io_out_d),
    .io_out_a(pCodeLock_io_out_a),
    .io_out_g(pCodeLock_io_out_g),
    .io_out_u(pCodeLock_io_out_u),
    .io_out_x(pCodeLock_io_out_x),
    .io_out_w(pCodeLock_io_out_w),
    .io_out_r(pCodeLock_io_out_r),
    .io_out_v(pCodeLock_io_out_v),
    .io_cfg_0_base(pCodeLock_io_cfg_0_base),
    .io_cfg_0_mask(pCodeLock_io_cfg_0_mask),
    .io_cfg_0_valid(pCodeLock_io_cfg_0_valid),
    .io_cfg_0_enable(pCodeLock_io_cfg_0_enable),
    .io_cfg_1_base(pCodeLock_io_cfg_1_base),
    .io_cfg_1_mask(pCodeLock_io_cfg_1_mask),
    .io_cfg_1_valid(pCodeLock_io_cfg_1_valid),
    .io_cfg_1_enable(pCodeLock_io_cfg_1_enable),
    .io_cfg_2_base(pCodeLock_io_cfg_2_base),
    .io_cfg_2_mask(pCodeLock_io_cfg_2_mask),
    .io_cfg_2_valid(pCodeLock_io_cfg_2_valid),
    .io_cfg_2_enable(pCodeLock_io_cfg_2_enable),
    .io_cfg_3_base(pCodeLock_io_cfg_3_base),
    .io_cfg_3_mask(pCodeLock_io_cfg_3_mask),
    .io_cfg_3_valid(pCodeLock_io_cfg_3_valid),
    .io_cfg_3_enable(pCodeLock_io_cfg_3_enable),
    .io_covSum(pCodeLock_io_covSum),
    .metaAssert(pCodeLock_metaAssert)
  );
  assign _T_582 = state != 3'h0; // @[PTW.scala 202:24]
  assign tmp_v = io_mem_resp_bits_data_word_bypass[0]; // @[PTW.scala 218:33]
  assign tmp_r = io_mem_resp_bits_data_word_bypass[1]; // @[PTW.scala 218:33]
  assign tmp_w = io_mem_resp_bits_data_word_bypass[2]; // @[PTW.scala 218:33]
  assign tmp_x = io_mem_resp_bits_data_word_bypass[3]; // @[PTW.scala 218:33]
  assign tmp_u = io_mem_resp_bits_data_word_bypass[4]; // @[PTW.scala 218:33]
  assign tmp_g = io_mem_resp_bits_data_word_bypass[5]; // @[PTW.scala 218:33]
  assign tmp_a = io_mem_resp_bits_data_word_bypass[6]; // @[PTW.scala 218:33]
  assign tmp_d = io_mem_resp_bits_data_word_bypass[7]; // @[PTW.scala 218:33]
  assign tmp_reserved_for_software = io_mem_resp_bits_data_word_bypass[9:8]; // @[PTW.scala 218:33]
  assign tmp_ppn = io_mem_resp_bits_data_word_bypass[63:10]; // @[PTW.scala 218:33]
  assign _T_624 = tmp_r | tmp_w; // @[PTW.scala 221:17]
  assign _T_625 = _T_624 | tmp_x; // @[PTW.scala 221:26]
  assign _T_626 = count <= 2'h0; // @[PTW.scala 224:21]
  assign _T_628 = tmp_ppn[17:9] != 9'h0; // @[PTW.scala 224:95]
  assign _T_629 = _T_626 & _T_628; // @[PTW.scala 224:26]
  assign _GEN_37 = _T_629 ? 1'h0 : tmp_v; // @[PTW.scala 224:102]
  assign _T_630 = count <= 2'h1; // @[PTW.scala 224:21]
  assign _T_632 = tmp_ppn[8:0] != 9'h0; // @[PTW.scala 224:95]
  assign _T_633 = _T_630 & _T_632; // @[PTW.scala 224:26]
  assign _GEN_38 = _T_633 ? 1'h0 : _GEN_37; // @[PTW.scala 224:102]
  assign res_v = _T_625 ? _GEN_38 : tmp_v; // @[PTW.scala 221:36]
  assign invalid_paddr = tmp_ppn[53:20] != 34'h0; // @[PTW.scala 226:32]
  assign _T_636 = res_v & ~tmp_r; // @[PTW.scala 76:33]
  assign _T_638 = _T_636 & ~tmp_w; // @[PTW.scala 76:39]
  assign _T_640 = _T_638 & ~tmp_x; // @[PTW.scala 76:45]
  assign _T_642 = _T_640 & ~invalid_paddr; // @[PTW.scala 228:30]
  assign _T_643 = count < 2'h2; // @[PTW.scala 228:57]
  assign traverse = _T_642 & _T_643; // @[PTW.scala 228:48]
  assign _T_650 = count == 2'h1; // @[package.scala 31:81]
  assign _T_651 = _T_650 ? r_req_addr[17:9] : r_req_addr[26:18]; // @[package.scala 31:71]
  assign _T_652 = count == 2'h2; // @[package.scala 31:81]
  assign _T_653 = _T_652 ? r_req_addr[8:0] : _T_651; // @[package.scala 31:71]
  assign _T_654 = count == 2'h3; // @[package.scala 31:81]
  assign vpn_idx = _T_654 ? r_req_addr[8:0] : _T_653; // @[package.scala 31:71]
  assign _T_655 = {r_pte_ppn,vpn_idx}; // @[Cat.scala 30:58]
  assign pte_addr = {_T_655, 3'h0}; // @[PTW.scala 232:29]
  assign _T_658 = {r_pte_ppn[53:6],r_req_addr[5:0]}; // @[Cat.scala 30:58]
  assign _T_661 = {r_pte_ppn[53:3],r_req_addr[2:0]}; // @[Cat.scala 30:58]
  assign fragmented_superpage_ppn = count[0] ? _T_661 : _T_658; // @[package.scala 31:71]
  assign _T_665 = arb_io_out_ready & arb_io_out_valid; // @[Decoupled.scala 37:37]
  assign valid = invalid ? 8'h0 : reg_valid; // @[PTW.scala 249:20]
  assign _GEN_148 = {{34'd0}, tags_0}; // @[PTW.scala 253:27]
  assign _T_696 = _GEN_148 == pte_addr; // @[PTW.scala 253:27]
  assign _GEN_149 = {{34'd0}, tags_1}; // @[PTW.scala 253:27]
  assign _T_697 = _GEN_149 == pte_addr; // @[PTW.scala 253:27]
  assign _GEN_150 = {{34'd0}, tags_2}; // @[PTW.scala 253:27]
  assign _T_698 = _GEN_150 == pte_addr; // @[PTW.scala 253:27]
  assign _GEN_151 = {{34'd0}, tags_3}; // @[PTW.scala 253:27]
  assign _T_699 = _GEN_151 == pte_addr; // @[PTW.scala 253:27]
  assign _GEN_152 = {{34'd0}, tags_4}; // @[PTW.scala 253:27]
  assign _T_700 = _GEN_152 == pte_addr; // @[PTW.scala 253:27]
  assign _GEN_153 = {{34'd0}, tags_5}; // @[PTW.scala 253:27]
  assign _T_701 = _GEN_153 == pte_addr; // @[PTW.scala 253:27]
  assign _GEN_154 = {{34'd0}, tags_6}; // @[PTW.scala 253:27]
  assign _T_702 = _GEN_154 == pte_addr; // @[PTW.scala 253:27]
  assign _GEN_155 = {{34'd0}, tags_7}; // @[PTW.scala 253:27]
  assign _T_703 = _GEN_155 == pte_addr; // @[PTW.scala 253:27]
  assign _T_710 = {_T_703,_T_702,_T_701,_T_700,_T_699,_T_698,_T_697,_T_696}; // @[Cat.scala 30:58]
  assign hits = _T_710 & valid; // @[PTW.scala 253:48]
  assign hit = hits != 8'h0; // @[PTW.scala 254:20]
  assign _T_711 = state == 3'h4; // @[PTW.scala 255:18]
  assign _T_712 = state == 3'h5; // @[PTW.scala 255:39]
  assign _T_713 = _T_711 | _T_712; // @[PTW.scala 255:30]
  assign _T_714 = _T_713 & traverse; // @[PTW.scala 255:52]
  assign _T_716 = _T_714 & ~hit; // @[PTW.scala 255:64]
  assign _T_718 = _T_716 & ~invalidated; // @[PTW.scala 255:72]
  assign _T_720 = ~valid == 8'h0; // @[PTW.scala 256:25]
  assign _T_721 = {_T_667, 1'h0}; // @[Replacement.scala 57:31]
  assign _T_725 = {{1'd0}, _T_721[7:1]}; // @[Replacement.scala 61:48]
  assign _T_728 = {1'h1,_T_725[0]}; // @[Cat.scala 30:58]
  assign _T_732 = _T_721 >> _T_728; // @[Replacement.scala 61:48]
  assign _T_735 = {1'h1,_T_725[0],_T_732[0]}; // @[Cat.scala 30:58]
  assign _T_739 = _T_721 >> _T_735; // @[Replacement.scala 61:48]
  assign _T_742 = {1'h1,_T_725[0],_T_732[0],_T_739[0]}; // @[Cat.scala 30:58]
  assign _T_745 = ~valid[0]; // @[OneHot.scala 39:40]
  assign _T_746 = ~valid[1]; // @[OneHot.scala 39:40]
  assign _T_747 = ~valid[2]; // @[OneHot.scala 39:40]
  assign _T_748 = ~valid[3]; // @[OneHot.scala 39:40]
  assign _T_749 = ~valid[4]; // @[OneHot.scala 39:40]
  assign _T_750 = ~valid[5]; // @[OneHot.scala 39:40]
  assign _T_751 = ~valid[6]; // @[OneHot.scala 39:40]
  assign _T_753 = _T_751 ? 3'h6 : 3'h7; // @[Mux.scala 31:69]
  assign _T_754 = _T_750 ? 3'h5 : _T_753; // @[Mux.scala 31:69]
  assign _T_755 = _T_749 ? 3'h4 : _T_754; // @[Mux.scala 31:69]
  assign _T_756 = _T_748 ? 3'h3 : _T_755; // @[Mux.scala 31:69]
  assign _T_757 = _T_747 ? 3'h2 : _T_756; // @[Mux.scala 31:69]
  assign _T_758 = _T_746 ? 3'h1 : _T_757; // @[Mux.scala 31:69]
  assign _T_759 = _T_745 ? 3'h0 : _T_758; // @[Mux.scala 31:69]
  assign r = _T_720 ? _T_742[2:0] : _T_759; // @[PTW.scala 256:18]
  assign _T_760 = 8'h1 << r; // @[OneHot.scala 45:35]
  assign _T_761 = valid | _T_760; // @[PTW.scala 258:49]
  assign _T_764 = valid & ~_T_760; // @[PTW.scala 258:70]
  assign res_ppn = {{34'd0}, tmp_ppn[19:0]}; // @[PTW.scala 220:13]
  assign _GEN_58 = _T_718 ? 1'h0 : invalid; // @[PTW.scala 255:89]
  assign _T_768 = state == 3'h1; // @[PTW.scala 262:24]
  assign _T_769 = hit & _T_768; // @[PTW.scala 262:15]
  assign _T_772 = hits[7:4] != 4'h0; // @[OneHot.scala 28:14]
  assign _T_773 = hits[7:4] | hits[3:0]; // @[OneHot.scala 28:28]
  assign _T_776 = _T_773[3:2] != 2'h0; // @[OneHot.scala 28:14]
  assign _T_777 = _T_773[3:2] | _T_773[1:0]; // @[OneHot.scala 28:28]
  assign _T_780 = {_T_772,_T_776,_T_777[1]}; // @[Cat.scala 30:58]
  assign _T_785 = _T_721 | 8'h2; // @[Replacement.scala 50:37]
  assign _T_787 = ~_T_721 | 8'h2; // @[Replacement.scala 50:37]
  assign _T_789 = _T_780[2] ? ~_T_787 : _T_785; // @[Replacement.scala 50:37]
  assign _T_790 = {1'h1,_T_780[2]}; // @[Cat.scala 30:58]
  assign _T_793 = 4'h1 << _T_790; // @[Replacement.scala 50:37]
  assign _GEN_157 = {{4'd0}, _T_793}; // @[Replacement.scala 50:37]
  assign _T_794 = _T_789 | _GEN_157; // @[Replacement.scala 50:37]
  assign _T_796 = ~_T_789 | _GEN_157; // @[Replacement.scala 50:37]
  assign _T_798 = _T_780[1] ? ~_T_796 : _T_794; // @[Replacement.scala 50:37]
  assign _T_799 = {1'h1,_T_780[2],_T_780[1]}; // @[Cat.scala 30:58]
  assign _T_802 = 8'h1 << _T_799; // @[Replacement.scala 50:37]
  assign _T_803 = _T_798 | _T_802; // @[Replacement.scala 50:37]
  assign _T_805 = ~_T_798 | _T_802; // @[Replacement.scala 50:37]
  assign _T_807 = _T_780[0] ? ~_T_805 : _T_803; // @[Replacement.scala 50:37]
  assign _T_811 = io_dpath_sfence_valid & ~io_dpath_sfence_bits_rs1; // @[PTW.scala 263:33]
  assign _GEN_77 = _T_811 | _GEN_58; // @[PTW.scala 263:63]
  assign pte_cache_hit = hit & _T_643; // @[PTW.scala 268:10]
  assign _T_830 = hits[0] ? data_0 : 20'h0; // @[Mux.scala 19:72]
  assign _T_831 = hits[1] ? data_1 : 20'h0; // @[Mux.scala 19:72]
  assign _T_832 = hits[2] ? data_2 : 20'h0; // @[Mux.scala 19:72]
  assign _T_833 = hits[3] ? data_3 : 20'h0; // @[Mux.scala 19:72]
  assign _T_834 = hits[4] ? data_4 : 20'h0; // @[Mux.scala 19:72]
  assign _T_835 = hits[5] ? data_5 : 20'h0; // @[Mux.scala 19:72]
  assign _T_836 = hits[6] ? data_6 : 20'h0; // @[Mux.scala 19:72]
  assign _T_837 = hits[7] ? data_7 : 20'h0; // @[Mux.scala 19:72]
  assign _T_838 = _T_830 | _T_831; // @[Mux.scala 19:72]
  assign _T_839 = _T_838 | _T_832; // @[Mux.scala 19:72]
  assign _T_840 = _T_839 | _T_833; // @[Mux.scala 19:72]
  assign _T_841 = _T_840 | _T_834; // @[Mux.scala 19:72]
  assign _T_842 = _T_841 | _T_835; // @[Mux.scala 19:72]
  assign _T_843 = _T_842 | _T_836; // @[Mux.scala 19:72]
  assign pte_cache_data = _T_843 | _T_837; // @[Mux.scala 19:72]
  assign _T_849 = invalidated & _T_582; // @[PTW.scala 341:56]
  assign _T_852 = state == 3'h3; // @[PTW.scala 343:48]
  assign _T_862 = pte_addr ^ 66'h60000000; // @[Parameters.scala 121:31]
  assign _T_863 = {1'b0,$signed(_T_862)}; // @[Parameters.scala 121:49]
  assign _T_865 = $signed(_T_863) & -67'sh20000000; // @[Parameters.scala 121:52]
  assign _T_866 = $signed(_T_865) == 67'sh0; // @[Parameters.scala 121:67]
  assign _T_867 = pte_addr ^ 66'hc000000; // @[Parameters.scala 121:31]
  assign _T_868 = {1'b0,$signed(_T_867)}; // @[Parameters.scala 121:49]
  assign _T_870 = $signed(_T_868) & -67'sh4000000; // @[Parameters.scala 121:52]
  assign _T_871 = $signed(_T_870) == 67'sh0; // @[Parameters.scala 121:67]
  assign _T_872 = pte_addr ^ 66'h80000000; // @[Parameters.scala 121:31]
  assign _T_873 = {1'b0,$signed(_T_872)}; // @[Parameters.scala 121:49]
  assign _T_875 = $signed(_T_873) & -67'sh10000000; // @[Parameters.scala 121:52]
  assign _T_876 = $signed(_T_875) == 67'sh0; // @[Parameters.scala 121:67]
  assign _T_878 = _T_866 | _T_871; // @[TLBPermissions.scala 97:65]
  assign _T_879 = _T_878 | _T_876; // @[TLBPermissions.scala 97:65]
  assign _T_883 = {1'b0,$signed(pte_addr)}; // @[Parameters.scala 121:49]
  assign _T_912 = pte_addr ^ 66'h3000; // @[Parameters.scala 121:31]
  assign _T_913 = {1'b0,$signed(_T_912)}; // @[Parameters.scala 121:49]
  assign _T_915 = $signed(_T_913) & -67'sh1000; // @[Parameters.scala 121:52]
  assign _T_916 = $signed(_T_915) == 67'sh0; // @[Parameters.scala 121:67]
  assign _T_922 = pte_addr ^ 66'h2000000; // @[Parameters.scala 121:31]
  assign _T_923 = {1'b0,$signed(_T_922)}; // @[Parameters.scala 121:49]
  assign _T_925 = $signed(_T_923) & -67'sh10000; // @[Parameters.scala 121:52]
  assign _T_926 = $signed(_T_925) == 67'sh0; // @[Parameters.scala 121:67]
  assign _T_927 = pte_addr ^ 66'h10000; // @[Parameters.scala 121:31]
  assign _T_928 = {1'b0,$signed(_T_927)}; // @[Parameters.scala 121:49]
  assign _T_930 = $signed(_T_928) & -67'sh10000; // @[Parameters.scala 121:52]
  assign _T_931 = $signed(_T_930) == 67'sh0; // @[Parameters.scala 121:67]
  assign _T_940 = $signed(_T_883) & -67'sh1000; // @[Parameters.scala 121:52]
  assign _T_941 = $signed(_T_940) == 67'sh0; // @[Parameters.scala 121:67]
  assign _T_943 = _T_866 | _T_916; // @[TLBPermissions.scala 97:65]
  assign _T_944 = _T_943 | _T_871; // @[TLBPermissions.scala 97:65]
  assign _T_945 = _T_944 | _T_926; // @[TLBPermissions.scala 97:65]
  assign _T_946 = _T_945 | _T_931; // @[TLBPermissions.scala 97:65]
  assign _T_947 = _T_946 | _T_876; // @[TLBPermissions.scala 97:65]
  assign _T_948 = _T_947 | _T_941; // @[TLBPermissions.scala 97:65]
  assign _T_1001 = _T_650 & _T_879; // @[package.scala 31:71]
  assign _T_1003 = _T_652 ? _T_948 : _T_1001; // @[package.scala 31:71]
  assign pmaHomogeneous = _T_654 ? _T_948 : _T_1003; // @[package.scala 31:71]
  assign _T_1006 = {pte_addr[65:12], 12'h0}; // @[PTW.scala 362:92]
  assign _T_1025 = _T_650 ? io_dpath_pmp_0_mask[20] : io_dpath_pmp_0_mask[29]; // @[package.scala 31:71]
  assign _T_1027 = _T_652 ? io_dpath_pmp_0_mask[11] : _T_1025; // @[package.scala 31:71]
  assign _T_1029 = _T_654 ? io_dpath_pmp_0_mask[11] : _T_1027; // @[package.scala 31:71]
  assign _T_1030 = {io_dpath_pmp_0_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_1032 = ~_T_1030 | 32'h3; // @[PMP.scala 54:48]
  assign _GEN_159 = {{34'd0}, ~_T_1032}; // @[PMP.scala 92:53]
  assign _T_1034 = _T_1006 ^ _GEN_159; // @[PMP.scala 92:53]
  assign _T_1036 = _T_1034[65:30] != 36'h0; // @[PMP.scala 92:78]
  assign _T_1043 = _T_1034[65:21] != 45'h0; // @[PMP.scala 92:78]
  assign _T_1050 = _T_1034[65:12] != 54'h0; // @[PMP.scala 92:78]
  assign _T_1052 = _T_650 ? _T_1043 : _T_1036; // @[package.scala 31:71]
  assign _T_1054 = _T_652 ? _T_1050 : _T_1052; // @[package.scala 31:71]
  assign _T_1056 = _T_654 ? _T_1050 : _T_1054; // @[package.scala 31:71]
  assign _T_1057 = _T_1029 | _T_1056; // @[PMP.scala 92:21]
  assign _T_1070 = _T_1006 < _GEN_159; // @[PMP.scala 101:32]
  assign _T_1073 = _T_650 ? 32'hffe00000 : 32'hc0000000; // @[package.scala 31:71]
  assign _T_1075 = _T_652 ? 32'hfffff000 : _T_1073; // @[package.scala 31:71]
  assign _T_1077 = _T_654 ? 32'hfffff000 : _T_1075; // @[package.scala 31:71]
  assign _GEN_163 = {{34'd0}, _T_1077}; // @[PMP.scala 104:30]
  assign _T_1078 = _T_1006 & _GEN_163; // @[PMP.scala 104:30]
  assign _T_1090 = ~_T_1032 & _T_1077; // @[PMP.scala 105:53]
  assign _GEN_165 = {{34'd0}, _T_1090}; // @[PMP.scala 105:40]
  assign _T_1091 = _T_1078 < _GEN_165; // @[PMP.scala 105:40]
  assign _T_1094 = ~_T_1070 | _T_1091; // @[PMP.scala 107:41]
  assign _T_1095 = ~io_dpath_pmp_0_cfg_a[0] | _T_1094; // @[PMP.scala 112:58]
  assign _T_1096 = io_dpath_pmp_0_cfg_a[1] ? _T_1057 : _T_1095; // @[PMP.scala 112:8]
  assign _T_1103 = _T_650 ? io_dpath_pmp_1_mask[20] : io_dpath_pmp_1_mask[29]; // @[package.scala 31:71]
  assign _T_1105 = _T_652 ? io_dpath_pmp_1_mask[11] : _T_1103; // @[package.scala 31:71]
  assign _T_1107 = _T_654 ? io_dpath_pmp_1_mask[11] : _T_1105; // @[package.scala 31:71]
  assign _T_1108 = {io_dpath_pmp_1_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_1110 = ~_T_1108 | 32'h3; // @[PMP.scala 54:48]
  assign _GEN_166 = {{34'd0}, ~_T_1110}; // @[PMP.scala 92:53]
  assign _T_1112 = _T_1006 ^ _GEN_166; // @[PMP.scala 92:53]
  assign _T_1114 = _T_1112[65:30] != 36'h0; // @[PMP.scala 92:78]
  assign _T_1121 = _T_1112[65:21] != 45'h0; // @[PMP.scala 92:78]
  assign _T_1128 = _T_1112[65:12] != 54'h0; // @[PMP.scala 92:78]
  assign _T_1130 = _T_650 ? _T_1121 : _T_1114; // @[package.scala 31:71]
  assign _T_1132 = _T_652 ? _T_1128 : _T_1130; // @[package.scala 31:71]
  assign _T_1134 = _T_654 ? _T_1128 : _T_1132; // @[package.scala 31:71]
  assign _T_1135 = _T_1107 | _T_1134; // @[PMP.scala 92:21]
  assign _T_1148 = _T_1006 < _GEN_166; // @[PMP.scala 101:32]
  assign _T_1168 = ~_T_1110 & _T_1077; // @[PMP.scala 105:53]
  assign _GEN_174 = {{34'd0}, _T_1168}; // @[PMP.scala 105:40]
  assign _T_1169 = _T_1078 < _GEN_174; // @[PMP.scala 105:40]
  assign _T_1170 = _T_1091 | ~_T_1148; // @[PMP.scala 107:21]
  assign _T_1171 = ~_T_1070 & _T_1169; // @[PMP.scala 107:62]
  assign _T_1172 = _T_1170 | _T_1171; // @[PMP.scala 107:41]
  assign _T_1173 = ~io_dpath_pmp_1_cfg_a[0] | _T_1172; // @[PMP.scala 112:58]
  assign _T_1174 = io_dpath_pmp_1_cfg_a[1] ? _T_1135 : _T_1173; // @[PMP.scala 112:8]
  assign _T_1175 = _T_1096 & _T_1174; // @[PMP.scala 132:10]
  assign _T_1181 = _T_650 ? io_dpath_pmp_2_mask[20] : io_dpath_pmp_2_mask[29]; // @[package.scala 31:71]
  assign _T_1183 = _T_652 ? io_dpath_pmp_2_mask[11] : _T_1181; // @[package.scala 31:71]
  assign _T_1185 = _T_654 ? io_dpath_pmp_2_mask[11] : _T_1183; // @[package.scala 31:71]
  assign _T_1186 = {io_dpath_pmp_2_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_1188 = ~_T_1186 | 32'h3; // @[PMP.scala 54:48]
  assign _GEN_175 = {{34'd0}, ~_T_1188}; // @[PMP.scala 92:53]
  assign _T_1190 = _T_1006 ^ _GEN_175; // @[PMP.scala 92:53]
  assign _T_1192 = _T_1190[65:30] != 36'h0; // @[PMP.scala 92:78]
  assign _T_1199 = _T_1190[65:21] != 45'h0; // @[PMP.scala 92:78]
  assign _T_1206 = _T_1190[65:12] != 54'h0; // @[PMP.scala 92:78]
  assign _T_1208 = _T_650 ? _T_1199 : _T_1192; // @[package.scala 31:71]
  assign _T_1210 = _T_652 ? _T_1206 : _T_1208; // @[package.scala 31:71]
  assign _T_1212 = _T_654 ? _T_1206 : _T_1210; // @[package.scala 31:71]
  assign _T_1213 = _T_1185 | _T_1212; // @[PMP.scala 92:21]
  assign _T_1226 = _T_1006 < _GEN_175; // @[PMP.scala 101:32]
  assign _T_1246 = ~_T_1188 & _T_1077; // @[PMP.scala 105:53]
  assign _GEN_183 = {{34'd0}, _T_1246}; // @[PMP.scala 105:40]
  assign _T_1247 = _T_1078 < _GEN_183; // @[PMP.scala 105:40]
  assign _T_1248 = _T_1169 | ~_T_1226; // @[PMP.scala 107:21]
  assign _T_1249 = ~_T_1148 & _T_1247; // @[PMP.scala 107:62]
  assign _T_1250 = _T_1248 | _T_1249; // @[PMP.scala 107:41]
  assign _T_1251 = ~io_dpath_pmp_2_cfg_a[0] | _T_1250; // @[PMP.scala 112:58]
  assign _T_1252 = io_dpath_pmp_2_cfg_a[1] ? _T_1213 : _T_1251; // @[PMP.scala 112:8]
  assign _T_1253 = _T_1175 & _T_1252; // @[PMP.scala 132:10]
  assign _T_1259 = _T_650 ? io_dpath_pmp_3_mask[20] : io_dpath_pmp_3_mask[29]; // @[package.scala 31:71]
  assign _T_1261 = _T_652 ? io_dpath_pmp_3_mask[11] : _T_1259; // @[package.scala 31:71]
  assign _T_1263 = _T_654 ? io_dpath_pmp_3_mask[11] : _T_1261; // @[package.scala 31:71]
  assign _T_1264 = {io_dpath_pmp_3_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_1266 = ~_T_1264 | 32'h3; // @[PMP.scala 54:48]
  assign _GEN_184 = {{34'd0}, ~_T_1266}; // @[PMP.scala 92:53]
  assign _T_1268 = _T_1006 ^ _GEN_184; // @[PMP.scala 92:53]
  assign _T_1270 = _T_1268[65:30] != 36'h0; // @[PMP.scala 92:78]
  assign _T_1277 = _T_1268[65:21] != 45'h0; // @[PMP.scala 92:78]
  assign _T_1284 = _T_1268[65:12] != 54'h0; // @[PMP.scala 92:78]
  assign _T_1286 = _T_650 ? _T_1277 : _T_1270; // @[package.scala 31:71]
  assign _T_1288 = _T_652 ? _T_1284 : _T_1286; // @[package.scala 31:71]
  assign _T_1290 = _T_654 ? _T_1284 : _T_1288; // @[package.scala 31:71]
  assign _T_1291 = _T_1263 | _T_1290; // @[PMP.scala 92:21]
  assign _T_1304 = _T_1006 < _GEN_184; // @[PMP.scala 101:32]
  assign _T_1324 = ~_T_1266 & _T_1077; // @[PMP.scala 105:53]
  assign _GEN_192 = {{34'd0}, _T_1324}; // @[PMP.scala 105:40]
  assign _T_1325 = _T_1078 < _GEN_192; // @[PMP.scala 105:40]
  assign _T_1326 = _T_1247 | ~_T_1304; // @[PMP.scala 107:21]
  assign _T_1327 = ~_T_1226 & _T_1325; // @[PMP.scala 107:62]
  assign _T_1328 = _T_1326 | _T_1327; // @[PMP.scala 107:41]
  assign _T_1329 = ~io_dpath_pmp_3_cfg_a[0] | _T_1328; // @[PMP.scala 112:58]
  assign _T_1330 = io_dpath_pmp_3_cfg_a[1] ? _T_1291 : _T_1329; // @[PMP.scala 112:8]
  assign _T_1331 = _T_1253 & _T_1330; // @[PMP.scala 132:10]
  assign _T_1337 = _T_650 ? io_dpath_pmp_4_mask[20] : io_dpath_pmp_4_mask[29]; // @[package.scala 31:71]
  assign _T_1339 = _T_652 ? io_dpath_pmp_4_mask[11] : _T_1337; // @[package.scala 31:71]
  assign _T_1341 = _T_654 ? io_dpath_pmp_4_mask[11] : _T_1339; // @[package.scala 31:71]
  assign _T_1342 = {io_dpath_pmp_4_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_1344 = ~_T_1342 | 32'h3; // @[PMP.scala 54:48]
  assign _GEN_193 = {{34'd0}, ~_T_1344}; // @[PMP.scala 92:53]
  assign _T_1346 = _T_1006 ^ _GEN_193; // @[PMP.scala 92:53]
  assign _T_1348 = _T_1346[65:30] != 36'h0; // @[PMP.scala 92:78]
  assign _T_1355 = _T_1346[65:21] != 45'h0; // @[PMP.scala 92:78]
  assign _T_1362 = _T_1346[65:12] != 54'h0; // @[PMP.scala 92:78]
  assign _T_1364 = _T_650 ? _T_1355 : _T_1348; // @[package.scala 31:71]
  assign _T_1366 = _T_652 ? _T_1362 : _T_1364; // @[package.scala 31:71]
  assign _T_1368 = _T_654 ? _T_1362 : _T_1366; // @[package.scala 31:71]
  assign _T_1369 = _T_1341 | _T_1368; // @[PMP.scala 92:21]
  assign _T_1382 = _T_1006 < _GEN_193; // @[PMP.scala 101:32]
  assign _T_1402 = ~_T_1344 & _T_1077; // @[PMP.scala 105:53]
  assign _GEN_201 = {{34'd0}, _T_1402}; // @[PMP.scala 105:40]
  assign _T_1403 = _T_1078 < _GEN_201; // @[PMP.scala 105:40]
  assign _T_1404 = _T_1325 | ~_T_1382; // @[PMP.scala 107:21]
  assign _T_1405 = ~_T_1304 & _T_1403; // @[PMP.scala 107:62]
  assign _T_1406 = _T_1404 | _T_1405; // @[PMP.scala 107:41]
  assign _T_1407 = ~io_dpath_pmp_4_cfg_a[0] | _T_1406; // @[PMP.scala 112:58]
  assign _T_1408 = io_dpath_pmp_4_cfg_a[1] ? _T_1369 : _T_1407; // @[PMP.scala 112:8]
  assign _T_1409 = _T_1331 & _T_1408; // @[PMP.scala 132:10]
  assign _T_1415 = _T_650 ? io_dpath_pmp_5_mask[20] : io_dpath_pmp_5_mask[29]; // @[package.scala 31:71]
  assign _T_1417 = _T_652 ? io_dpath_pmp_5_mask[11] : _T_1415; // @[package.scala 31:71]
  assign _T_1419 = _T_654 ? io_dpath_pmp_5_mask[11] : _T_1417; // @[package.scala 31:71]
  assign _T_1420 = {io_dpath_pmp_5_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_1422 = ~_T_1420 | 32'h3; // @[PMP.scala 54:48]
  assign _GEN_202 = {{34'd0}, ~_T_1422}; // @[PMP.scala 92:53]
  assign _T_1424 = _T_1006 ^ _GEN_202; // @[PMP.scala 92:53]
  assign _T_1426 = _T_1424[65:30] != 36'h0; // @[PMP.scala 92:78]
  assign _T_1433 = _T_1424[65:21] != 45'h0; // @[PMP.scala 92:78]
  assign _T_1440 = _T_1424[65:12] != 54'h0; // @[PMP.scala 92:78]
  assign _T_1442 = _T_650 ? _T_1433 : _T_1426; // @[package.scala 31:71]
  assign _T_1444 = _T_652 ? _T_1440 : _T_1442; // @[package.scala 31:71]
  assign _T_1446 = _T_654 ? _T_1440 : _T_1444; // @[package.scala 31:71]
  assign _T_1447 = _T_1419 | _T_1446; // @[PMP.scala 92:21]
  assign _T_1460 = _T_1006 < _GEN_202; // @[PMP.scala 101:32]
  assign _T_1480 = ~_T_1422 & _T_1077; // @[PMP.scala 105:53]
  assign _GEN_210 = {{34'd0}, _T_1480}; // @[PMP.scala 105:40]
  assign _T_1481 = _T_1078 < _GEN_210; // @[PMP.scala 105:40]
  assign _T_1482 = _T_1403 | ~_T_1460; // @[PMP.scala 107:21]
  assign _T_1483 = ~_T_1382 & _T_1481; // @[PMP.scala 107:62]
  assign _T_1484 = _T_1482 | _T_1483; // @[PMP.scala 107:41]
  assign _T_1485 = ~io_dpath_pmp_5_cfg_a[0] | _T_1484; // @[PMP.scala 112:58]
  assign _T_1486 = io_dpath_pmp_5_cfg_a[1] ? _T_1447 : _T_1485; // @[PMP.scala 112:8]
  assign _T_1487 = _T_1409 & _T_1486; // @[PMP.scala 132:10]
  assign _T_1493 = _T_650 ? io_dpath_pmp_6_mask[20] : io_dpath_pmp_6_mask[29]; // @[package.scala 31:71]
  assign _T_1495 = _T_652 ? io_dpath_pmp_6_mask[11] : _T_1493; // @[package.scala 31:71]
  assign _T_1497 = _T_654 ? io_dpath_pmp_6_mask[11] : _T_1495; // @[package.scala 31:71]
  assign _T_1498 = {io_dpath_pmp_6_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_1500 = ~_T_1498 | 32'h3; // @[PMP.scala 54:48]
  assign _GEN_211 = {{34'd0}, ~_T_1500}; // @[PMP.scala 92:53]
  assign _T_1502 = _T_1006 ^ _GEN_211; // @[PMP.scala 92:53]
  assign _T_1504 = _T_1502[65:30] != 36'h0; // @[PMP.scala 92:78]
  assign _T_1511 = _T_1502[65:21] != 45'h0; // @[PMP.scala 92:78]
  assign _T_1518 = _T_1502[65:12] != 54'h0; // @[PMP.scala 92:78]
  assign _T_1520 = _T_650 ? _T_1511 : _T_1504; // @[package.scala 31:71]
  assign _T_1522 = _T_652 ? _T_1518 : _T_1520; // @[package.scala 31:71]
  assign _T_1524 = _T_654 ? _T_1518 : _T_1522; // @[package.scala 31:71]
  assign _T_1525 = _T_1497 | _T_1524; // @[PMP.scala 92:21]
  assign _T_1538 = _T_1006 < _GEN_211; // @[PMP.scala 101:32]
  assign _T_1558 = ~_T_1500 & _T_1077; // @[PMP.scala 105:53]
  assign _GEN_219 = {{34'd0}, _T_1558}; // @[PMP.scala 105:40]
  assign _T_1559 = _T_1078 < _GEN_219; // @[PMP.scala 105:40]
  assign _T_1560 = _T_1481 | ~_T_1538; // @[PMP.scala 107:21]
  assign _T_1561 = ~_T_1460 & _T_1559; // @[PMP.scala 107:62]
  assign _T_1562 = _T_1560 | _T_1561; // @[PMP.scala 107:41]
  assign _T_1563 = ~io_dpath_pmp_6_cfg_a[0] | _T_1562; // @[PMP.scala 112:58]
  assign _T_1564 = io_dpath_pmp_6_cfg_a[1] ? _T_1525 : _T_1563; // @[PMP.scala 112:8]
  assign _T_1565 = _T_1487 & _T_1564; // @[PMP.scala 132:10]
  assign _T_1571 = _T_650 ? io_dpath_pmp_7_mask[20] : io_dpath_pmp_7_mask[29]; // @[package.scala 31:71]
  assign _T_1573 = _T_652 ? io_dpath_pmp_7_mask[11] : _T_1571; // @[package.scala 31:71]
  assign _T_1575 = _T_654 ? io_dpath_pmp_7_mask[11] : _T_1573; // @[package.scala 31:71]
  assign _T_1576 = {io_dpath_pmp_7_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_1578 = ~_T_1576 | 32'h3; // @[PMP.scala 54:48]
  assign _GEN_220 = {{34'd0}, ~_T_1578}; // @[PMP.scala 92:53]
  assign _T_1580 = _T_1006 ^ _GEN_220; // @[PMP.scala 92:53]
  assign _T_1582 = _T_1580[65:30] != 36'h0; // @[PMP.scala 92:78]
  assign _T_1589 = _T_1580[65:21] != 45'h0; // @[PMP.scala 92:78]
  assign _T_1596 = _T_1580[65:12] != 54'h0; // @[PMP.scala 92:78]
  assign _T_1598 = _T_650 ? _T_1589 : _T_1582; // @[package.scala 31:71]
  assign _T_1600 = _T_652 ? _T_1596 : _T_1598; // @[package.scala 31:71]
  assign _T_1602 = _T_654 ? _T_1596 : _T_1600; // @[package.scala 31:71]
  assign _T_1603 = _T_1575 | _T_1602; // @[PMP.scala 92:21]
  assign _T_1616 = _T_1006 < _GEN_220; // @[PMP.scala 101:32]
  assign _T_1636 = ~_T_1578 & _T_1077; // @[PMP.scala 105:53]
  assign _GEN_228 = {{34'd0}, _T_1636}; // @[PMP.scala 105:40]
  assign _T_1637 = _T_1078 < _GEN_228; // @[PMP.scala 105:40]
  assign _T_1638 = _T_1559 | ~_T_1616; // @[PMP.scala 107:21]
  assign _T_1639 = ~_T_1538 & _T_1637; // @[PMP.scala 107:62]
  assign _T_1640 = _T_1638 | _T_1639; // @[PMP.scala 107:41]
  assign _T_1641 = ~io_dpath_pmp_7_cfg_a[0] | _T_1640; // @[PMP.scala 112:58]
  assign _T_1642 = io_dpath_pmp_7_cfg_a[1] ? _T_1603 : _T_1641; // @[PMP.scala 112:8]
  assign pmpHomogeneous = _T_1565 & _T_1642; // @[PMP.scala 132:10]
  assign homogeneous = pmaHomogeneous & pmpHomogeneous; // @[PTW.scala 363:36]
  assign ae = res_v & invalid_paddr; // @[PTW.scala 492:22]
  assign _GEN_136 = traverse ? 3'h1 : 3'h0; // @[PTW.scala 487:21]
  assign _T_1650 = 3'h0 == state; // @[Conditional.scala 37:30]
  assign _T_1652 = arb_io_out_bits_valid ? 3'h1 : 3'h0; // @[PTW.scala 393:26]
  assign _GEN_80 = _T_665 ? _T_1652 : state; // @[PTW.scala 392:32]
  assign _T_1653 = 3'h1 == state; // @[Conditional.scala 37:30]
  assign _T_1656 = io_mem_req_ready ? 3'h2 : 3'h1; // @[PTW.scala 401:26]
  assign _GEN_82 = pte_cache_hit ? state : _T_1656; // @[PTW.scala 398:28]
  assign _T_1657 = 3'h2 == state; // @[Conditional.scala 37:30]
  assign _T_1658 = 3'h4 == state; // @[Conditional.scala 37:30]
  assign _GEN_86 = io_mem_s2_xcpt_ae_ld ? 3'h0 : 3'h5; // @[PTW.scala 409:35]
  assign _T_1664 = 3'h7 == state; // @[Conditional.scala 37:30]
  assign _GEN_93 = _T_1664 ? 3'h0 : state; // @[Conditional.scala 39:67]
  assign _GEN_99 = _T_1658 ? _GEN_86 : _GEN_93; // @[Conditional.scala 39:67]
  assign _GEN_105 = _T_1657 ? 3'h4 : _GEN_99; // @[Conditional.scala 39:67]
  assign _GEN_112 = _T_1653 ? _GEN_82 : _GEN_105; // @[Conditional.scala 39:67]
  assign _GEN_117 = _T_1650 ? _GEN_80 : _GEN_112; // @[Conditional.scala 40:58]
  assign _GEN_130 = io_mem_s2_nack ? 3'h1 : _GEN_117; // @[PTW.scala 481:25]
  assign next_state = io_mem_resp_valid ? _GEN_136 : _GEN_130; // @[PTW.scala 485:28]
  assign _T_1655 = count + 2'h1; // @[PTW.scala 399:24]
  assign _GEN_87 = io_mem_s2_xcpt_ae_ld & ~r_req_dest; // @[PTW.scala 409:35]
  assign _GEN_88 = io_mem_s2_xcpt_ae_ld & r_req_dest; // @[PTW.scala 409:35]
  assign _GEN_94 = _T_1664 & ~r_req_dest; // @[Conditional.scala 39:67]
  assign _GEN_95 = _T_1664 & r_req_dest; // @[Conditional.scala 39:67]
  assign _GEN_100 = _T_1658 & io_mem_s2_xcpt_ae_ld; // @[Conditional.scala 39:67]
  assign _GEN_101 = _T_1658 ? _GEN_87 : _GEN_94; // @[Conditional.scala 39:67]
  assign _GEN_102 = _T_1658 ? _GEN_88 : _GEN_95; // @[Conditional.scala 39:67]
  assign _GEN_107 = _T_1657 ? 1'h0 : _GEN_101; // @[Conditional.scala 39:67]
  assign _GEN_108 = _T_1657 ? 1'h0 : _GEN_102; // @[Conditional.scala 39:67]
  assign _GEN_114 = _T_1653 ? 1'h0 : _GEN_107; // @[Conditional.scala 39:67]
  assign _GEN_115 = _T_1653 ? 1'h0 : _GEN_108; // @[Conditional.scala 39:67]
  assign _GEN_120 = _T_1650 ? 1'h0 : _GEN_114; // @[Conditional.scala 40:58]
  assign _GEN_121 = _T_1650 ? 1'h0 : _GEN_115; // @[Conditional.scala 40:58]
  assign _T_1671 = state == 3'h7; // @[PTW.scala 465:15]
  assign _T_1673 = _T_1671 & ~homogeneous; // @[PTW.scala 465:40]
  assign _T_1676 = _T_768 & pte_cache_hit; // @[PTW.scala 466:25]
  assign pte_2_ppn = {{10'd0}, io_dpath_ptbr_ppn}; // @[PTW.scala 428:13]
  assign _T_1680_ppn = _T_665 ? pte_2_ppn : r_pte_ppn; // @[PTW.scala 467:8]
  assign pte_1_ppn = {{34'd0}, pte_cache_data}; // @[PTW.scala 428:13]
  assign _T_1681_ppn = _T_1676 ? pte_1_ppn : _T_1680_ppn; // @[PTW.scala 466:8]
  assign _T_1681_reserved_for_software = _T_1676 ? 2'h0 : r_pte_reserved_for_software; // @[PTW.scala 466:8]
  assign _T_1681_d = _T_1676 ? 1'h0 : r_pte_d; // @[PTW.scala 466:8]
  assign _T_1681_a = _T_1676 ? 1'h0 : r_pte_a; // @[PTW.scala 466:8]
  assign _T_1681_g = _T_1676 ? 1'h0 : r_pte_g; // @[PTW.scala 466:8]
  assign _T_1681_u = _T_1676 ? 1'h0 : r_pte_u; // @[PTW.scala 466:8]
  assign _T_1681_x = _T_1676 ? 1'h0 : r_pte_x; // @[PTW.scala 466:8]
  assign _T_1681_w = _T_1676 ? 1'h0 : r_pte_w; // @[PTW.scala 466:8]
  assign _T_1681_r = _T_1676 ? 1'h0 : r_pte_r; // @[PTW.scala 466:8]
  assign _T_1681_v = _T_1676 ? 1'h0 : r_pte_v; // @[PTW.scala 466:8]
  assign _T_1682_ppn = _T_1673 ? fragmented_superpage_ppn : _T_1681_ppn; // @[PTW.scala 465:8]
  assign _T_1682_reserved_for_software = _T_1673 ? r_pte_reserved_for_software : _T_1681_reserved_for_software; // @[PTW.scala 465:8]
  assign _T_1682_d = _T_1673 ? r_pte_d : _T_1681_d; // @[PTW.scala 465:8]
  assign _T_1682_a = _T_1673 ? r_pte_a : _T_1681_a; // @[PTW.scala 465:8]
  assign _T_1682_g = _T_1673 ? r_pte_g : _T_1681_g; // @[PTW.scala 465:8]
  assign _T_1682_u = _T_1673 ? r_pte_u : _T_1681_u; // @[PTW.scala 465:8]
  assign _T_1682_x = _T_1673 ? r_pte_x : _T_1681_x; // @[PTW.scala 465:8]
  assign _T_1682_w = _T_1673 ? r_pte_w : _T_1681_w; // @[PTW.scala 465:8]
  assign _T_1682_r = _T_1673 ? r_pte_r : _T_1681_r; // @[PTW.scala 465:8]
  assign _T_1682_v = _T_1673 ? r_pte_v : _T_1681_v; // @[PTW.scala 465:8]
  assign _T_1684_ppn = io_mem_resp_valid ? res_ppn : _T_1682_ppn; // @[PTW.scala 463:8]
  assign _T_1684_reserved_for_software = io_mem_resp_valid ? tmp_reserved_for_software : _T_1682_reserved_for_software; // @[PTW.scala 463:8]
  assign _T_1684_d = io_mem_resp_valid ? tmp_d : _T_1682_d; // @[PTW.scala 463:8]
  assign _T_1684_a = io_mem_resp_valid ? tmp_a : _T_1682_a; // @[PTW.scala 463:8]
  assign _T_1684_g = io_mem_resp_valid ? tmp_g : _T_1682_g; // @[PTW.scala 463:8]
  assign _T_1684_u = io_mem_resp_valid ? tmp_u : _T_1682_u; // @[PTW.scala 463:8]
  assign _T_1684_x = io_mem_resp_valid ? tmp_x : _T_1682_x; // @[PTW.scala 463:8]
  assign _T_1684_w = io_mem_resp_valid ? tmp_w : _T_1682_w; // @[PTW.scala 463:8]
  assign _T_1684_r = io_mem_resp_valid ? tmp_r : _T_1682_r; // @[PTW.scala 463:8]
  assign _T_1684_v = io_mem_resp_valid ? res_v : _T_1682_v; // @[PTW.scala 463:8]
  assign _T_1693 = {_T_1684_ppn,_T_1684_reserved_for_software,_T_1684_d,_T_1684_a,_T_1684_g,_T_1684_u,_T_1684_x,_T_1684_w,_T_1684_r,_T_1684_v}; // @[package.scala 208:71]
  assign _GEN_123 = ~r_req_dest | _GEN_120; // @[PTW.scala 477:28]
  assign _GEN_124 = r_req_dest | _GEN_121; // @[PTW.scala 477:28]
  assign _T_1723 = _T_711 | reset; // @[PTW.scala 482:11]
  assign _T_1729 = _T_713 | reset; // @[PTW.scala 486:11]
  assign io_requestor_0_req_ready = arb_io_in_0_ready; // @[PTW.scala 198:13]
  assign io_requestor_0_resp_valid = resp_valid_0; // @[PTW.scala 374:32]
  assign io_requestor_0_resp_bits_ae = resp_ae; // @[PTW.scala 375:34]
  assign io_requestor_0_resp_bits_pte_ppn = r_pte_ppn; // @[PTW.scala 376:35]
  assign io_requestor_0_resp_bits_pte_d = r_pte_d; // @[PTW.scala 376:35]
  assign io_requestor_0_resp_bits_pte_a = r_pte_a; // @[PTW.scala 376:35]
  assign io_requestor_0_resp_bits_pte_g = r_pte_g; // @[PTW.scala 376:35]
  assign io_requestor_0_resp_bits_pte_u = r_pte_u; // @[PTW.scala 376:35]
  assign io_requestor_0_resp_bits_pte_x = r_pte_x; // @[PTW.scala 376:35]
  assign io_requestor_0_resp_bits_pte_w = r_pte_w; // @[PTW.scala 376:35]
  assign io_requestor_0_resp_bits_pte_r = r_pte_r; // @[PTW.scala 376:35]
  assign io_requestor_0_resp_bits_pte_v = r_pte_v; // @[PTW.scala 376:35]
  assign io_requestor_0_resp_bits_level = count; // @[PTW.scala 377:37]
  assign io_requestor_0_resp_bits_homogeneous = pmaHomogeneous & pmpHomogeneous; // @[PTW.scala 378:43]
  assign io_requestor_0_ptbr_mode = io_dpath_ptbr_mode; // @[PTW.scala 380:26]
  assign io_requestor_0_status_dprv = io_dpath_status_dprv; // @[PTW.scala 382:28]
  assign io_requestor_0_status_mxr = io_dpath_status_mxr; // @[PTW.scala 382:28]
  assign io_requestor_0_status_sum = io_dpath_status_sum; // @[PTW.scala 382:28]
  assign io_requestor_0_pmp_0_cfg_l = io_dpath_pmp_0_cfg_l; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_0_cfg_a = io_dpath_pmp_0_cfg_a; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_0_cfg_x = io_dpath_pmp_0_cfg_x; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_0_cfg_w = io_dpath_pmp_0_cfg_w; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_0_cfg_r = io_dpath_pmp_0_cfg_r; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_0_addr = io_dpath_pmp_0_addr; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_0_mask = io_dpath_pmp_0_mask; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_1_cfg_l = io_dpath_pmp_1_cfg_l; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_1_cfg_a = io_dpath_pmp_1_cfg_a; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_1_cfg_x = io_dpath_pmp_1_cfg_x; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_1_cfg_w = io_dpath_pmp_1_cfg_w; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_1_cfg_r = io_dpath_pmp_1_cfg_r; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_1_addr = io_dpath_pmp_1_addr; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_1_mask = io_dpath_pmp_1_mask; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_2_cfg_l = io_dpath_pmp_2_cfg_l; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_2_cfg_a = io_dpath_pmp_2_cfg_a; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_2_cfg_x = io_dpath_pmp_2_cfg_x; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_2_cfg_w = io_dpath_pmp_2_cfg_w; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_2_cfg_r = io_dpath_pmp_2_cfg_r; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_2_addr = io_dpath_pmp_2_addr; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_2_mask = io_dpath_pmp_2_mask; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_3_cfg_l = io_dpath_pmp_3_cfg_l; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_3_cfg_a = io_dpath_pmp_3_cfg_a; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_3_cfg_x = io_dpath_pmp_3_cfg_x; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_3_cfg_w = io_dpath_pmp_3_cfg_w; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_3_cfg_r = io_dpath_pmp_3_cfg_r; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_3_addr = io_dpath_pmp_3_addr; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_3_mask = io_dpath_pmp_3_mask; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_4_cfg_l = io_dpath_pmp_4_cfg_l; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_4_cfg_a = io_dpath_pmp_4_cfg_a; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_4_cfg_x = io_dpath_pmp_4_cfg_x; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_4_cfg_w = io_dpath_pmp_4_cfg_w; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_4_cfg_r = io_dpath_pmp_4_cfg_r; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_4_addr = io_dpath_pmp_4_addr; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_4_mask = io_dpath_pmp_4_mask; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_5_cfg_l = io_dpath_pmp_5_cfg_l; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_5_cfg_a = io_dpath_pmp_5_cfg_a; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_5_cfg_x = io_dpath_pmp_5_cfg_x; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_5_cfg_w = io_dpath_pmp_5_cfg_w; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_5_cfg_r = io_dpath_pmp_5_cfg_r; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_5_addr = io_dpath_pmp_5_addr; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_5_mask = io_dpath_pmp_5_mask; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_6_cfg_l = io_dpath_pmp_6_cfg_l; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_6_cfg_a = io_dpath_pmp_6_cfg_a; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_6_cfg_x = io_dpath_pmp_6_cfg_x; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_6_cfg_w = io_dpath_pmp_6_cfg_w; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_6_cfg_r = io_dpath_pmp_6_cfg_r; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_6_addr = io_dpath_pmp_6_addr; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_6_mask = io_dpath_pmp_6_mask; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_7_cfg_l = io_dpath_pmp_7_cfg_l; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_7_cfg_a = io_dpath_pmp_7_cfg_a; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_7_cfg_x = io_dpath_pmp_7_cfg_x; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_7_cfg_w = io_dpath_pmp_7_cfg_w; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_7_cfg_r = io_dpath_pmp_7_cfg_r; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_7_addr = io_dpath_pmp_7_addr; // @[PTW.scala 383:25]
  assign io_requestor_0_pmp_7_mask = io_dpath_pmp_7_mask; // @[PTW.scala 383:25]
  assign io_requestor_0_vpoffset_bits_value = io_dpath_vpoffset_req_bits_value; // @[PTW.scala 370:45]
  assign io_requestor_1_req_ready = arb_io_in_1_ready; // @[PTW.scala 198:13]
  assign io_requestor_1_resp_valid = resp_valid_1; // @[PTW.scala 374:32]
  assign io_requestor_1_resp_bits_ae = resp_ae; // @[PTW.scala 375:34]
  assign io_requestor_1_resp_bits_pte_ppn = r_pte_ppn; // @[PTW.scala 376:35]
  assign io_requestor_1_resp_bits_pte_d = r_pte_d; // @[PTW.scala 376:35]
  assign io_requestor_1_resp_bits_pte_a = r_pte_a; // @[PTW.scala 376:35]
  assign io_requestor_1_resp_bits_pte_g = r_pte_g; // @[PTW.scala 376:35]
  assign io_requestor_1_resp_bits_pte_u = r_pte_u; // @[PTW.scala 376:35]
  assign io_requestor_1_resp_bits_pte_x = r_pte_x; // @[PTW.scala 376:35]
  assign io_requestor_1_resp_bits_pte_w = r_pte_w; // @[PTW.scala 376:35]
  assign io_requestor_1_resp_bits_pte_r = r_pte_r; // @[PTW.scala 376:35]
  assign io_requestor_1_resp_bits_pte_v = r_pte_v; // @[PTW.scala 376:35]
  assign io_requestor_1_resp_bits_level = count; // @[PTW.scala 377:37]
  assign io_requestor_1_resp_bits_homogeneous = pmaHomogeneous & pmpHomogeneous; // @[PTW.scala 378:43]
  assign io_requestor_1_ptbr_mode = io_dpath_ptbr_mode; // @[PTW.scala 380:26]
  assign io_requestor_1_status_prv = io_dpath_status_prv; // @[PTW.scala 382:28]
  assign io_requestor_1_pmp_0_cfg_l = io_dpath_pmp_0_cfg_l; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_0_cfg_a = io_dpath_pmp_0_cfg_a; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_0_cfg_x = io_dpath_pmp_0_cfg_x; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_0_cfg_w = io_dpath_pmp_0_cfg_w; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_0_cfg_r = io_dpath_pmp_0_cfg_r; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_0_addr = io_dpath_pmp_0_addr; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_0_mask = io_dpath_pmp_0_mask; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_1_cfg_l = io_dpath_pmp_1_cfg_l; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_1_cfg_a = io_dpath_pmp_1_cfg_a; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_1_cfg_x = io_dpath_pmp_1_cfg_x; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_1_cfg_w = io_dpath_pmp_1_cfg_w; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_1_cfg_r = io_dpath_pmp_1_cfg_r; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_1_addr = io_dpath_pmp_1_addr; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_1_mask = io_dpath_pmp_1_mask; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_2_cfg_l = io_dpath_pmp_2_cfg_l; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_2_cfg_a = io_dpath_pmp_2_cfg_a; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_2_cfg_x = io_dpath_pmp_2_cfg_x; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_2_cfg_w = io_dpath_pmp_2_cfg_w; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_2_cfg_r = io_dpath_pmp_2_cfg_r; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_2_addr = io_dpath_pmp_2_addr; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_2_mask = io_dpath_pmp_2_mask; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_3_cfg_l = io_dpath_pmp_3_cfg_l; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_3_cfg_a = io_dpath_pmp_3_cfg_a; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_3_cfg_x = io_dpath_pmp_3_cfg_x; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_3_cfg_w = io_dpath_pmp_3_cfg_w; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_3_cfg_r = io_dpath_pmp_3_cfg_r; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_3_addr = io_dpath_pmp_3_addr; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_3_mask = io_dpath_pmp_3_mask; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_4_cfg_l = io_dpath_pmp_4_cfg_l; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_4_cfg_a = io_dpath_pmp_4_cfg_a; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_4_cfg_x = io_dpath_pmp_4_cfg_x; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_4_cfg_w = io_dpath_pmp_4_cfg_w; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_4_cfg_r = io_dpath_pmp_4_cfg_r; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_4_addr = io_dpath_pmp_4_addr; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_4_mask = io_dpath_pmp_4_mask; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_5_cfg_l = io_dpath_pmp_5_cfg_l; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_5_cfg_a = io_dpath_pmp_5_cfg_a; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_5_cfg_x = io_dpath_pmp_5_cfg_x; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_5_cfg_w = io_dpath_pmp_5_cfg_w; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_5_cfg_r = io_dpath_pmp_5_cfg_r; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_5_addr = io_dpath_pmp_5_addr; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_5_mask = io_dpath_pmp_5_mask; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_6_cfg_l = io_dpath_pmp_6_cfg_l; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_6_cfg_a = io_dpath_pmp_6_cfg_a; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_6_cfg_x = io_dpath_pmp_6_cfg_x; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_6_cfg_w = io_dpath_pmp_6_cfg_w; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_6_cfg_r = io_dpath_pmp_6_cfg_r; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_6_addr = io_dpath_pmp_6_addr; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_6_mask = io_dpath_pmp_6_mask; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_7_cfg_l = io_dpath_pmp_7_cfg_l; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_7_cfg_a = io_dpath_pmp_7_cfg_a; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_7_cfg_x = io_dpath_pmp_7_cfg_x; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_7_cfg_w = io_dpath_pmp_7_cfg_w; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_7_cfg_r = io_dpath_pmp_7_cfg_r; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_7_addr = io_dpath_pmp_7_addr; // @[PTW.scala 383:25]
  assign io_requestor_1_pmp_7_mask = io_dpath_pmp_7_mask; // @[PTW.scala 383:25]
  assign io_requestor_1_vpoffset_bits_value = io_dpath_vpoffset_req_bits_value; // @[PTW.scala 370:45]
  assign io_mem_req_valid = _T_768 | _T_852; // @[PTW.scala 343:20]
  assign io_mem_req_bits_addr = pte_addr[39:0]; // @[PTW.scala 347:24]
  assign io_mem_s1_kill = state != 3'h2; // @[PTW.scala 348:18]
  assign arb_clock = clock;
  assign arb_io_in_0_valid = io_requestor_0_req_valid; // @[PTW.scala 198:13]
  assign arb_io_in_0_bits_bits_addr = io_requestor_0_req_bits_bits_addr; // @[PTW.scala 198:13]
  assign arb_io_in_1_valid = io_requestor_1_req_valid; // @[PTW.scala 198:13]
  assign arb_io_in_1_bits_valid = io_requestor_1_req_bits_valid; // @[PTW.scala 198:13]
  assign arb_io_in_1_bits_bits_addr = io_requestor_1_req_bits_bits_addr; // @[PTW.scala 198:13]
  assign arb_io_out_ready = state == 3'h0; // @[PTW.scala 199:20]
  assign pCodeLock_io_in_ppn = _T_1693[63:10]; // @[PTW.scala 471:19]
  assign pCodeLock_io_in_reserved_for_software = _T_1693[9:8]; // @[PTW.scala 471:19]
  assign pCodeLock_io_in_d = _T_1693[7]; // @[PTW.scala 471:19]
  assign pCodeLock_io_in_a = _T_1693[6]; // @[PTW.scala 471:19]
  assign pCodeLock_io_in_g = _T_1693[5]; // @[PTW.scala 471:19]
  assign pCodeLock_io_in_u = _T_1693[4]; // @[PTW.scala 471:19]
  assign pCodeLock_io_in_x = _T_1693[3]; // @[PTW.scala 471:19]
  assign pCodeLock_io_in_w = _T_1693[2]; // @[PTW.scala 471:19]
  assign pCodeLock_io_in_r = _T_1693[1]; // @[PTW.scala 471:19]
  assign pCodeLock_io_in_v = _T_1693[0]; // @[PTW.scala 471:19]
  assign pCodeLock_io_cfg_0_base = pcode_cfg_0_base; // @[PTW.scala 470:20]
  assign pCodeLock_io_cfg_0_mask = pcode_cfg_0_mask; // @[PTW.scala 470:20]
  assign pCodeLock_io_cfg_0_valid = pcode_cfg_0_valid; // @[PTW.scala 470:20]
  assign pCodeLock_io_cfg_0_enable = pcode_cfg_0_enable; // @[PTW.scala 470:20]
  assign pCodeLock_io_cfg_1_base = pcode_cfg_1_base; // @[PTW.scala 470:20]
  assign pCodeLock_io_cfg_1_mask = pcode_cfg_1_mask; // @[PTW.scala 470:20]
  assign pCodeLock_io_cfg_1_valid = pcode_cfg_1_valid; // @[PTW.scala 470:20]
  assign pCodeLock_io_cfg_1_enable = pcode_cfg_1_enable; // @[PTW.scala 470:20]
  assign pCodeLock_io_cfg_2_base = pcode_cfg_2_base; // @[PTW.scala 470:20]
  assign pCodeLock_io_cfg_2_mask = pcode_cfg_2_mask; // @[PTW.scala 470:20]
  assign pCodeLock_io_cfg_2_valid = pcode_cfg_2_valid; // @[PTW.scala 470:20]
  assign pCodeLock_io_cfg_2_enable = pcode_cfg_2_enable; // @[PTW.scala 470:20]
  assign pCodeLock_io_cfg_3_base = pcode_cfg_3_base; // @[PTW.scala 470:20]
  assign pCodeLock_io_cfg_3_mask = pcode_cfg_3_mask; // @[PTW.scala 470:20]
  assign pCodeLock_io_cfg_3_valid = pcode_cfg_3_valid; // @[PTW.scala 470:20]
  assign pCodeLock_io_cfg_3_enable = pcode_cfg_3_enable; // @[PTW.scala 470:20]
  assign PTW_cov_read_addr = PTW_state;
  assign PTW_cov_read_data = PTW_cov[PTW_cov_read_addr]; // @[Coverage map for PTW]
  assign PTW_cov_write_data = 1'h1;
  assign PTW_cov_write_addr = PTW_state;
  assign PTW_cov_write_mask = 1'h1;
  assign PTW_cov_write_en = 1'h1;
  assign count_shl = {count, 15'h0};
  assign count_pad = {3'h0,count_shl};
  assign invalid_shl = {invalid, 10'h0};
  assign invalid_pad = {9'h0,invalid_shl};
  assign state_shl = {state, 8'h0};
  assign state_pad = {9'h0,state_shl};
  assign reg_valid_shl = {reg_valid, 2'h0};
  assign reg_valid_pad = {10'h0,reg_valid_shl};
  assign _T_667_shl = {_T_667, 3'h0};
  assign _T_667_pad = {10'h0,_T_667_shl};
  assign invalidated_shl = {invalidated, 8'h0};
  assign invalidated_pad = {11'h0,invalidated_shl};
  assign pcode_cfg_0_enable_shl = {pcode_cfg_0_enable, 12'h0};
  assign pcode_cfg_0_enable_pad = {7'h0,pcode_cfg_0_enable_shl};
  assign pcode_cfg_0_base_shl = pcode_cfg_0_base;
  assign pcode_cfg_0_base_pad = pcode_cfg_0_base_shl;
  assign pcode_cfg_0_mask_shl = {pcode_cfg_0_mask, 6'h0};
  assign pcode_cfg_0_mask_pad = {4'h0,pcode_cfg_0_mask_shl};
  assign pcode_cfg_0_valid_shl = {pcode_cfg_0_valid, 1'h0};
  assign pcode_cfg_0_valid_pad = {18'h0,pcode_cfg_0_valid_shl};
  assign PTW_xor3 = count_pad ^ invalid_pad;
  assign PTW_xor10 = reg_valid_pad ^ _T_667_pad;
  assign PTW_xor4 = state_pad ^ PTW_xor10;
  assign PTW_xor1 = PTW_xor3 ^ PTW_xor4;
  assign PTW_xor5 = invalidated_pad ^ pcode_cfg_0_enable_pad;
  assign PTW_xor14 = pcode_cfg_0_mask_pad ^ pcode_cfg_0_valid_pad;
  assign PTW_xor6 = pcode_cfg_0_base_pad ^ PTW_xor14;
  assign PTW_xor2 = PTW_xor5 ^ PTW_xor6;
  assign PTW_xor0 = PTW_xor1 ^ PTW_xor2;
  assign arb_sum = PTW_covSum + arb_io_covSum;
  assign pCodeLock_sum = arb_sum + pCodeLock_io_covSum;
  assign io_covSum = pCodeLock_sum;
  assign stopEn0 = io_mem_s2_nack & ~_T_1723;
  assign stopEn1 = io_mem_resp_valid & ~_T_1729;
  assign arb_metaAssert_wire = arb_metaAssert;
  assign pCodeLock_metaAssert_wire = pCodeLock_metaAssert;
  assign PTW_or1 = stopEn0 | stopEn1;
  assign PTW_or2 = arb_metaAssert_wire | pCodeLock_metaAssert_wire;
  assign PTW_or0 = PTW_or1 | PTW_or2;
  assign metaAssert = PTW_metaAssert;
  assign arb_metaReset = metaReset | arb_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pcode_cfg_0_base = _RAND_0[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  pcode_cfg_0_mask = _RAND_1[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  pcode_cfg_0_valid = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  pcode_cfg_0_enable = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  pcode_cfg_1_base = _RAND_4[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  pcode_cfg_1_mask = _RAND_5[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  pcode_cfg_1_valid = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  pcode_cfg_1_enable = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  pcode_cfg_2_base = _RAND_8[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  pcode_cfg_2_mask = _RAND_9[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  pcode_cfg_2_valid = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  pcode_cfg_2_enable = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  pcode_cfg_3_base = _RAND_12[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  pcode_cfg_3_mask = _RAND_13[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  pcode_cfg_3_valid = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  pcode_cfg_3_enable = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  state = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  resp_valid_0 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  resp_valid_1 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  invalidated = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  count = _RAND_20[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  resp_ae = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  r_req_addr = _RAND_22[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  r_req_dest = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {2{`RANDOM}};
  r_pte_ppn = _RAND_24[53:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  r_pte_reserved_for_software = _RAND_25[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  r_pte_d = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  r_pte_a = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  r_pte_g = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  r_pte_u = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  r_pte_x = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  r_pte_w = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  r_pte_r = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  r_pte_v = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_667 = _RAND_34[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  invalid = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  reg_valid = _RAND_36[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  tags_0 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  tags_1 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  tags_2 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  tags_3 = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  tags_4 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  tags_5 = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  tags_6 = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  tags_7 = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  data_0 = _RAND_45[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  data_1 = _RAND_46[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  data_2 = _RAND_47[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  data_3 = _RAND_48[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  data_4 = _RAND_49[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  data_5 = _RAND_50[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  data_6 = _RAND_51[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  data_7 = _RAND_52[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  PTW_state = _RAND_53[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    PTW_cov[initvar] = _RAND_54[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  PTW_covSum = _RAND_55[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  PTW_metaAssert = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      pcode_cfg_0_base <= 20'h0;
    end else if (reset) begin
      pcode_cfg_0_base <= 20'h0;
    end else if (io_dpath_pcode_req_valid) begin
      if (2'h0 == io_dpath_pcode_req_bits_id) begin
        pcode_cfg_0_base <= io_dpath_pcode_req_bits_value_base;
      end
    end
    if (metaReset) begin
      pcode_cfg_0_mask <= 10'h0;
    end else if (reset) begin
      pcode_cfg_0_mask <= 10'h0;
    end else if (io_dpath_pcode_req_valid) begin
      if (2'h0 == io_dpath_pcode_req_bits_id) begin
        pcode_cfg_0_mask <= io_dpath_pcode_req_bits_value_mask;
      end
    end
    if (metaReset) begin
      pcode_cfg_0_valid <= 1'h0;
    end else if (reset) begin
      pcode_cfg_0_valid <= 1'h0;
    end else if (io_dpath_pcode_req_valid) begin
      if (2'h0 == io_dpath_pcode_req_bits_id) begin
        pcode_cfg_0_valid <= io_dpath_pcode_req_bits_value_valid;
      end
    end
    if (metaReset) begin
      pcode_cfg_0_enable <= 1'h0;
    end else if (reset) begin
      pcode_cfg_0_enable <= 1'h0;
    end else if (io_dpath_pcode_req_valid) begin
      if (2'h0 == io_dpath_pcode_req_bits_id) begin
        pcode_cfg_0_enable <= io_dpath_pcode_req_bits_value_locked;
      end
    end
    if (metaReset) begin
      pcode_cfg_1_base <= 20'h0;
    end else if (reset) begin
      pcode_cfg_1_base <= 20'h0;
    end else if (io_dpath_pcode_req_valid) begin
      if (2'h1 == io_dpath_pcode_req_bits_id) begin
        pcode_cfg_1_base <= io_dpath_pcode_req_bits_value_base;
      end
    end
    if (metaReset) begin
      pcode_cfg_1_mask <= 10'h0;
    end else if (reset) begin
      pcode_cfg_1_mask <= 10'h0;
    end else if (io_dpath_pcode_req_valid) begin
      if (2'h1 == io_dpath_pcode_req_bits_id) begin
        pcode_cfg_1_mask <= io_dpath_pcode_req_bits_value_mask;
      end
    end
    if (metaReset) begin
      pcode_cfg_1_valid <= 1'h0;
    end else if (reset) begin
      pcode_cfg_1_valid <= 1'h0;
    end else if (io_dpath_pcode_req_valid) begin
      if (2'h1 == io_dpath_pcode_req_bits_id) begin
        pcode_cfg_1_valid <= io_dpath_pcode_req_bits_value_valid;
      end
    end
    if (metaReset) begin
      pcode_cfg_1_enable <= 1'h0;
    end else if (reset) begin
      pcode_cfg_1_enable <= 1'h0;
    end else if (io_dpath_pcode_req_valid) begin
      if (2'h1 == io_dpath_pcode_req_bits_id) begin
        pcode_cfg_1_enable <= io_dpath_pcode_req_bits_value_locked;
      end
    end
    if (metaReset) begin
      pcode_cfg_2_base <= 20'h0;
    end else if (reset) begin
      pcode_cfg_2_base <= 20'h0;
    end else if (io_dpath_pcode_req_valid) begin
      if (2'h2 == io_dpath_pcode_req_bits_id) begin
        pcode_cfg_2_base <= io_dpath_pcode_req_bits_value_base;
      end
    end
    if (metaReset) begin
      pcode_cfg_2_mask <= 10'h0;
    end else if (reset) begin
      pcode_cfg_2_mask <= 10'h0;
    end else if (io_dpath_pcode_req_valid) begin
      if (2'h2 == io_dpath_pcode_req_bits_id) begin
        pcode_cfg_2_mask <= io_dpath_pcode_req_bits_value_mask;
      end
    end
    if (metaReset) begin
      pcode_cfg_2_valid <= 1'h0;
    end else if (reset) begin
      pcode_cfg_2_valid <= 1'h0;
    end else if (io_dpath_pcode_req_valid) begin
      if (2'h2 == io_dpath_pcode_req_bits_id) begin
        pcode_cfg_2_valid <= io_dpath_pcode_req_bits_value_valid;
      end
    end
    if (metaReset) begin
      pcode_cfg_2_enable <= 1'h0;
    end else if (reset) begin
      pcode_cfg_2_enable <= 1'h0;
    end else if (io_dpath_pcode_req_valid) begin
      if (2'h2 == io_dpath_pcode_req_bits_id) begin
        pcode_cfg_2_enable <= io_dpath_pcode_req_bits_value_locked;
      end
    end
    if (metaReset) begin
      pcode_cfg_3_base <= 20'h0;
    end else if (reset) begin
      pcode_cfg_3_base <= 20'h0;
    end else if (io_dpath_pcode_req_valid) begin
      if (2'h3 == io_dpath_pcode_req_bits_id) begin
        pcode_cfg_3_base <= io_dpath_pcode_req_bits_value_base;
      end
    end
    if (metaReset) begin
      pcode_cfg_3_mask <= 10'h0;
    end else if (reset) begin
      pcode_cfg_3_mask <= 10'h0;
    end else if (io_dpath_pcode_req_valid) begin
      if (2'h3 == io_dpath_pcode_req_bits_id) begin
        pcode_cfg_3_mask <= io_dpath_pcode_req_bits_value_mask;
      end
    end
    if (metaReset) begin
      pcode_cfg_3_valid <= 1'h0;
    end else if (reset) begin
      pcode_cfg_3_valid <= 1'h0;
    end else if (io_dpath_pcode_req_valid) begin
      if (2'h3 == io_dpath_pcode_req_bits_id) begin
        pcode_cfg_3_valid <= io_dpath_pcode_req_bits_value_valid;
      end
    end
    if (metaReset) begin
      pcode_cfg_3_enable <= 1'h0;
    end else if (reset) begin
      pcode_cfg_3_enable <= 1'h0;
    end else if (io_dpath_pcode_req_valid) begin
      if (2'h3 == io_dpath_pcode_req_bits_id) begin
        pcode_cfg_3_enable <= io_dpath_pcode_req_bits_value_locked;
      end
    end
    if (metaReset) begin
      state <= 3'h0;
    end else if (reset) begin
      state <= 3'h0;
    end else begin
      state <= next_state[2:0];
    end
    if (metaReset) begin
      resp_valid_0 <= 1'h0;
    end else if (io_mem_resp_valid) begin
      if (traverse) begin
        if (_T_1650) begin
          resp_valid_0 <= 1'h0;
        end else if (_T_1653) begin
          resp_valid_0 <= 1'h0;
        end else if (_T_1657) begin
          resp_valid_0 <= 1'h0;
        end else if (_T_1658) begin
          resp_valid_0 <= _GEN_87;
        end else begin
          resp_valid_0 <= _GEN_94;
        end
      end else begin
        resp_valid_0 <= _GEN_123;
      end
    end else if (_T_1650) begin
      resp_valid_0 <= 1'h0;
    end else if (_T_1653) begin
      resp_valid_0 <= 1'h0;
    end else if (_T_1657) begin
      resp_valid_0 <= 1'h0;
    end else if (_T_1658) begin
      resp_valid_0 <= _GEN_87;
    end else begin
      resp_valid_0 <= _GEN_94;
    end
    if (metaReset) begin
      resp_valid_1 <= 1'h0;
    end else if (io_mem_resp_valid) begin
      if (traverse) begin
        if (_T_1650) begin
          resp_valid_1 <= 1'h0;
        end else if (_T_1653) begin
          resp_valid_1 <= 1'h0;
        end else if (_T_1657) begin
          resp_valid_1 <= 1'h0;
        end else if (_T_1658) begin
          resp_valid_1 <= _GEN_88;
        end else begin
          resp_valid_1 <= _GEN_95;
        end
      end else begin
        resp_valid_1 <= _GEN_124;
      end
    end else if (_T_1650) begin
      resp_valid_1 <= 1'h0;
    end else if (_T_1653) begin
      resp_valid_1 <= 1'h0;
    end else if (_T_1657) begin
      resp_valid_1 <= 1'h0;
    end else if (_T_1658) begin
      resp_valid_1 <= _GEN_88;
    end else begin
      resp_valid_1 <= _GEN_95;
    end
    if (metaReset) begin
      invalidated <= 1'h0;
    end else begin
      invalidated <= io_dpath_sfence_valid | _T_849;
    end
    if (metaReset) begin
      count <= 2'h0;
    end else if (io_mem_resp_valid) begin
      if (traverse) begin
        count <= _T_1655;
      end else if (_T_1650) begin
        count <= 2'h0;
      end else if (_T_1653) begin
        if (pte_cache_hit) begin
          count <= _T_1655;
        end
      end else if (!(_T_1657)) begin
        if (!(_T_1658)) begin
          if (_T_1664) begin
            if (~homogeneous) begin
              count <= 2'h2;
            end
          end
        end
      end
    end else if (_T_1650) begin
      count <= 2'h0;
    end else if (_T_1653) begin
      if (pte_cache_hit) begin
        count <= _T_1655;
      end
    end else if (!(_T_1657)) begin
      if (!(_T_1658)) begin
        if (_T_1664) begin
          if (~homogeneous) begin
            count <= 2'h2;
          end
        end
      end
    end
    if (metaReset) begin
      resp_ae <= 1'h0;
    end else if (io_mem_resp_valid) begin
      if (traverse) begin
        if (_T_1650) begin
          resp_ae <= 1'h0;
        end else if (_T_1653) begin
          resp_ae <= 1'h0;
        end else if (_T_1657) begin
          resp_ae <= 1'h0;
        end else begin
          resp_ae <= _GEN_100;
        end
      end else begin
        resp_ae <= ae;
      end
    end else if (_T_1650) begin
      resp_ae <= 1'h0;
    end else if (_T_1653) begin
      resp_ae <= 1'h0;
    end else if (_T_1657) begin
      resp_ae <= 1'h0;
    end else begin
      resp_ae <= _GEN_100;
    end
    if (metaReset) begin
      r_req_addr <= 27'h0;
    end else if (_T_665) begin
      r_req_addr <= arb_io_out_bits_bits_addr;
    end
    if (metaReset) begin
      r_req_dest <= 1'h0;
    end else if (_T_665) begin
      r_req_dest <= arb_io_chosen;
    end
    if (metaReset) begin
      r_pte_ppn <= 54'h0;
    end else begin
      r_pte_ppn <= pCodeLock_io_out_ppn;
    end
    if (metaReset) begin
      r_pte_reserved_for_software <= 2'h0;
    end else begin
      r_pte_reserved_for_software <= pCodeLock_io_out_reserved_for_software;
    end
    if (metaReset) begin
      r_pte_d <= 1'h0;
    end else begin
      r_pte_d <= pCodeLock_io_out_d;
    end
    if (metaReset) begin
      r_pte_a <= 1'h0;
    end else begin
      r_pte_a <= pCodeLock_io_out_a;
    end
    if (metaReset) begin
      r_pte_g <= 1'h0;
    end else begin
      r_pte_g <= pCodeLock_io_out_g;
    end
    if (metaReset) begin
      r_pte_u <= 1'h0;
    end else begin
      r_pte_u <= pCodeLock_io_out_u;
    end
    if (metaReset) begin
      r_pte_x <= 1'h0;
    end else begin
      r_pte_x <= pCodeLock_io_out_x;
    end
    if (metaReset) begin
      r_pte_w <= 1'h0;
    end else begin
      r_pte_w <= pCodeLock_io_out_w;
    end
    if (metaReset) begin
      r_pte_r <= 1'h0;
    end else begin
      r_pte_r <= pCodeLock_io_out_r;
    end
    if (metaReset) begin
      r_pte_v <= 1'h0;
    end else begin
      r_pte_v <= pCodeLock_io_out_v;
    end
    if (metaReset) begin
      _T_667 <= 7'h0;
    end else if (_T_769) begin
      _T_667 <= _T_807[7:1];
    end
    if (metaReset) begin
      invalid <= 1'h0;
    end else begin
      invalid <= reset | _GEN_77;
    end
    if (metaReset) begin
      reg_valid <= 8'h0;
    end else if (_T_718) begin
      if (io_mem_resp_valid) begin
        reg_valid <= _T_761;
      end else begin
        reg_valid <= _T_764;
      end
    end
    if (metaReset) begin
      tags_0 <= 32'h0;
    end else if (_T_718) begin
      if (3'h0 == r) begin
        tags_0 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      tags_1 <= 32'h0;
    end else if (_T_718) begin
      if (3'h1 == r) begin
        tags_1 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      tags_2 <= 32'h0;
    end else if (_T_718) begin
      if (3'h2 == r) begin
        tags_2 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      tags_3 <= 32'h0;
    end else if (_T_718) begin
      if (3'h3 == r) begin
        tags_3 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      tags_4 <= 32'h0;
    end else if (_T_718) begin
      if (3'h4 == r) begin
        tags_4 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      tags_5 <= 32'h0;
    end else if (_T_718) begin
      if (3'h5 == r) begin
        tags_5 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      tags_6 <= 32'h0;
    end else if (_T_718) begin
      if (3'h6 == r) begin
        tags_6 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      tags_7 <= 32'h0;
    end else if (_T_718) begin
      if (3'h7 == r) begin
        tags_7 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      data_0 <= 20'h0;
    end else if (_T_718) begin
      if (3'h0 == r) begin
        data_0 <= res_ppn[19:0];
      end
    end
    if (metaReset) begin
      data_1 <= 20'h0;
    end else if (_T_718) begin
      if (3'h1 == r) begin
        data_1 <= res_ppn[19:0];
      end
    end
    if (metaReset) begin
      data_2 <= 20'h0;
    end else if (_T_718) begin
      if (3'h2 == r) begin
        data_2 <= res_ppn[19:0];
      end
    end
    if (metaReset) begin
      data_3 <= 20'h0;
    end else if (_T_718) begin
      if (3'h3 == r) begin
        data_3 <= res_ppn[19:0];
      end
    end
    if (metaReset) begin
      data_4 <= 20'h0;
    end else if (_T_718) begin
      if (3'h4 == r) begin
        data_4 <= res_ppn[19:0];
      end
    end
    if (metaReset) begin
      data_5 <= 20'h0;
    end else if (_T_718) begin
      if (3'h5 == r) begin
        data_5 <= res_ppn[19:0];
      end
    end
    if (metaReset) begin
      data_6 <= 20'h0;
    end else if (_T_718) begin
      if (3'h6 == r) begin
        data_6 <= res_ppn[19:0];
      end
    end
    if (metaReset) begin
      data_7 <= 20'h0;
    end else if (_T_718) begin
      if (3'h7 == r) begin
        data_7 <= res_ppn[19:0];
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_mem_s2_nack & ~_T_1723) begin
          $fwrite(32'h80000002,"Assertion failed\n    at PTW.scala:482 assert(state === s_wait2)\n"); // @[PTW.scala 482:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_mem_s2_nack & ~_T_1723) begin
          $fatal; // @[PTW.scala 482:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_mem_resp_valid & ~_T_1729) begin
          $fwrite(32'h80000002,"Assertion failed\n    at PTW.scala:486 assert(state === s_wait2 || state === s_wait3)\n"); // @[PTW.scala 486:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_mem_resp_valid & ~_T_1729) begin
          $fatal; // @[PTW.scala 486:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    PTW_state <= PTW_xor0;
    if (!(PTW_cov_read_data)) begin
      PTW_covSum <= PTW_covSum + 1'h1;
    end
    if (metaReset) begin
      PTW_metaAssert <= 1'h0;
    end else begin
      PTW_metaAssert <= PTW_metaAssert | PTW_or0;
    end
  end
  always @(posedge clock) begin
    if(PTW_cov_write_en & PTW_cov_write_mask) begin
      PTW_cov[PTW_cov_write_addr] <= PTW_cov_write_data; // @[Coverage map for PTW]
    end
  end
endmodule
module Rocket(
  input         clock,
  input         reset,
  input  [1:0]  io_hartid,
  input         io_interrupts_debug,
  input         io_interrupts_mtip,
  input         io_interrupts_msip,
  input         io_interrupts_meip,
  input         io_interrupts_seip,
  output        io_imem_might_request,
  output        io_imem_req_valid,
  output [39:0] io_imem_req_bits_pc,
  output        io_imem_req_bits_speculative,
  output        io_imem_sfence_valid,
  output        io_imem_sfence_bits_rs1,
  output        io_imem_sfence_bits_rs2,
  output [38:0] io_imem_sfence_bits_addr,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input         io_imem_resp_bits_btb_taken,
  input         io_imem_resp_bits_btb_bridx,
  input  [4:0]  io_imem_resp_bits_btb_entry,
  input  [7:0]  io_imem_resp_bits_btb_bht_history,
  input  [39:0] io_imem_resp_bits_pc,
  input  [31:0] io_imem_resp_bits_data,
  input         io_imem_resp_bits_xcpt_pf_inst,
  input         io_imem_resp_bits_xcpt_ae_inst,
  input         io_imem_resp_bits_replay,
  output        io_imem_btb_update_valid,
  output [4:0]  io_imem_btb_update_bits_prediction_entry,
  output [38:0] io_imem_btb_update_bits_pc,
  output        io_imem_btb_update_bits_isValid,
  output [38:0] io_imem_btb_update_bits_br_pc,
  output [1:0]  io_imem_btb_update_bits_cfiType,
  output        io_imem_bht_update_valid,
  output [7:0]  io_imem_bht_update_bits_prediction_history,
  output [38:0] io_imem_bht_update_bits_pc,
  output        io_imem_bht_update_bits_branch,
  output        io_imem_bht_update_bits_taken,
  output        io_imem_bht_update_bits_mispredict,
  output        io_imem_flush_icache,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [39:0] io_dmem_req_bits_addr,
  output [6:0]  io_dmem_req_bits_tag,
  output [4:0]  io_dmem_req_bits_cmd,
  output [2:0]  io_dmem_req_bits_typ,
  output        io_dmem_s1_kill,
  output [63:0] io_dmem_s1_data_data,
  input         io_dmem_s2_nack,
  input         io_dmem_resp_valid,
  input  [6:0]  io_dmem_resp_bits_tag,
  input  [2:0]  io_dmem_resp_bits_typ,
  input  [63:0] io_dmem_resp_bits_data,
  input         io_dmem_resp_bits_replay,
  input         io_dmem_resp_bits_has_data,
  input  [63:0] io_dmem_resp_bits_data_word_bypass,
  input         io_dmem_replay_next,
  input         io_dmem_s2_xcpt_ma_ld,
  input         io_dmem_s2_xcpt_ma_st,
  input         io_dmem_s2_xcpt_pf_ld,
  input         io_dmem_s2_xcpt_pf_st,
  input         io_dmem_s2_xcpt_ae_ld,
  input         io_dmem_s2_xcpt_ae_st,
  input         io_dmem_ordered,
  input         io_dmem_perf_grant,
  output        io_dmem_keep_clock_enabled,
  input         io_dmem_clock_enabled,
  output [3:0]  io_ptw_ptbr_mode,
  output [43:0] io_ptw_ptbr_ppn,
  output        io_ptw_sfence_valid,
  output        io_ptw_sfence_bits_rs1,
  output [1:0]  io_ptw_status_dprv,
  output [1:0]  io_ptw_status_prv,
  output        io_ptw_status_mxr,
  output        io_ptw_status_sum,
  output        io_ptw_pmp_0_cfg_l,
  output [1:0]  io_ptw_pmp_0_cfg_a,
  output        io_ptw_pmp_0_cfg_x,
  output        io_ptw_pmp_0_cfg_w,
  output        io_ptw_pmp_0_cfg_r,
  output [29:0] io_ptw_pmp_0_addr,
  output [31:0] io_ptw_pmp_0_mask,
  output        io_ptw_pmp_1_cfg_l,
  output [1:0]  io_ptw_pmp_1_cfg_a,
  output        io_ptw_pmp_1_cfg_x,
  output        io_ptw_pmp_1_cfg_w,
  output        io_ptw_pmp_1_cfg_r,
  output [29:0] io_ptw_pmp_1_addr,
  output [31:0] io_ptw_pmp_1_mask,
  output        io_ptw_pmp_2_cfg_l,
  output [1:0]  io_ptw_pmp_2_cfg_a,
  output        io_ptw_pmp_2_cfg_x,
  output        io_ptw_pmp_2_cfg_w,
  output        io_ptw_pmp_2_cfg_r,
  output [29:0] io_ptw_pmp_2_addr,
  output [31:0] io_ptw_pmp_2_mask,
  output        io_ptw_pmp_3_cfg_l,
  output [1:0]  io_ptw_pmp_3_cfg_a,
  output        io_ptw_pmp_3_cfg_x,
  output        io_ptw_pmp_3_cfg_w,
  output        io_ptw_pmp_3_cfg_r,
  output [29:0] io_ptw_pmp_3_addr,
  output [31:0] io_ptw_pmp_3_mask,
  output        io_ptw_pmp_4_cfg_l,
  output [1:0]  io_ptw_pmp_4_cfg_a,
  output        io_ptw_pmp_4_cfg_x,
  output        io_ptw_pmp_4_cfg_w,
  output        io_ptw_pmp_4_cfg_r,
  output [29:0] io_ptw_pmp_4_addr,
  output [31:0] io_ptw_pmp_4_mask,
  output        io_ptw_pmp_5_cfg_l,
  output [1:0]  io_ptw_pmp_5_cfg_a,
  output        io_ptw_pmp_5_cfg_x,
  output        io_ptw_pmp_5_cfg_w,
  output        io_ptw_pmp_5_cfg_r,
  output [29:0] io_ptw_pmp_5_addr,
  output [31:0] io_ptw_pmp_5_mask,
  output        io_ptw_pmp_6_cfg_l,
  output [1:0]  io_ptw_pmp_6_cfg_a,
  output        io_ptw_pmp_6_cfg_x,
  output        io_ptw_pmp_6_cfg_w,
  output        io_ptw_pmp_6_cfg_r,
  output [29:0] io_ptw_pmp_6_addr,
  output [31:0] io_ptw_pmp_6_mask,
  output        io_ptw_pmp_7_cfg_l,
  output [1:0]  io_ptw_pmp_7_cfg_a,
  output        io_ptw_pmp_7_cfg_x,
  output        io_ptw_pmp_7_cfg_w,
  output        io_ptw_pmp_7_cfg_r,
  output [29:0] io_ptw_pmp_7_addr,
  output [31:0] io_ptw_pmp_7_mask,
  output [63:0] io_ptw_customCSRs_csrs_0_value,
  output        io_ptw_pcode_req_valid,
  output [1:0]  io_ptw_pcode_req_bits_id,
  output [19:0] io_ptw_pcode_req_bits_value_base,
  output [9:0]  io_ptw_pcode_req_bits_value_mask,
  output        io_ptw_pcode_req_bits_value_valid,
  output        io_ptw_pcode_req_bits_value_locked,
  output [26:0] io_ptw_vpoffset_req_bits_value,
  output [31:0] io_fpu_inst,
  output [63:0] io_fpu_fromint_data,
  output [2:0]  io_fpu_fcsr_rm,
  input         io_fpu_fcsr_flags_valid,
  input  [4:0]  io_fpu_fcsr_flags_bits,
  input  [63:0] io_fpu_store_data,
  input  [63:0] io_fpu_toint_data,
  output        io_fpu_dmem_resp_val,
  output [2:0]  io_fpu_dmem_resp_type,
  output [4:0]  io_fpu_dmem_resp_tag,
  output [63:0] io_fpu_dmem_resp_data,
  output        io_fpu_valid,
  input         io_fpu_fcsr_rdy,
  input         io_fpu_nack_mem,
  input         io_fpu_illegal_rm,
  output        io_fpu_killx,
  output        io_fpu_killm,
  input         io_fpu_dec_wen,
  input         io_fpu_dec_ren1,
  input         io_fpu_dec_ren2,
  input         io_fpu_dec_ren3,
  input         io_fpu_sboard_set,
  input         io_fpu_sboard_clr,
  input  [4:0]  io_fpu_sboard_clra,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         csr_halt,
  input         div_halt,
  input         ibuf_halt
);
  wire  ibuf_clock; // @[RocketCore.scala 236:20]
  wire  ibuf_reset; // @[RocketCore.scala 236:20]
  wire  ibuf_io_imem_ready; // @[RocketCore.scala 236:20]
  wire  ibuf_io_imem_valid; // @[RocketCore.scala 236:20]
  wire  ibuf_io_imem_bits_btb_taken; // @[RocketCore.scala 236:20]
  wire  ibuf_io_imem_bits_btb_bridx; // @[RocketCore.scala 236:20]
  wire [4:0] ibuf_io_imem_bits_btb_entry; // @[RocketCore.scala 236:20]
  wire [7:0] ibuf_io_imem_bits_btb_bht_history; // @[RocketCore.scala 236:20]
  wire [39:0] ibuf_io_imem_bits_pc; // @[RocketCore.scala 236:20]
  wire [31:0] ibuf_io_imem_bits_data; // @[RocketCore.scala 236:20]
  wire  ibuf_io_imem_bits_xcpt_pf_inst; // @[RocketCore.scala 236:20]
  wire  ibuf_io_imem_bits_xcpt_ae_inst; // @[RocketCore.scala 236:20]
  wire  ibuf_io_imem_bits_replay; // @[RocketCore.scala 236:20]
  wire  ibuf_io_kill; // @[RocketCore.scala 236:20]
  wire [39:0] ibuf_io_pc; // @[RocketCore.scala 236:20]
  wire [4:0] ibuf_io_btb_resp_entry; // @[RocketCore.scala 236:20]
  wire [7:0] ibuf_io_btb_resp_bht_history; // @[RocketCore.scala 236:20]
  wire  ibuf_io_inst_0_ready; // @[RocketCore.scala 236:20]
  wire  ibuf_io_inst_0_valid; // @[RocketCore.scala 236:20]
  wire  ibuf_io_inst_0_bits_xcpt0_pf_inst; // @[RocketCore.scala 236:20]
  wire  ibuf_io_inst_0_bits_xcpt0_ae_inst; // @[RocketCore.scala 236:20]
  wire  ibuf_io_inst_0_bits_xcpt1_pf_inst; // @[RocketCore.scala 236:20]
  wire  ibuf_io_inst_0_bits_xcpt1_ae_inst; // @[RocketCore.scala 236:20]
  wire  ibuf_io_inst_0_bits_replay; // @[RocketCore.scala 236:20]
  wire  ibuf_io_inst_0_bits_rvc; // @[RocketCore.scala 236:20]
  wire [31:0] ibuf_io_inst_0_bits_inst_bits; // @[RocketCore.scala 236:20]
  wire [4:0] ibuf_io_inst_0_bits_inst_rd; // @[RocketCore.scala 236:20]
  wire [4:0] ibuf_io_inst_0_bits_inst_rs1; // @[RocketCore.scala 236:20]
  wire [4:0] ibuf_io_inst_0_bits_inst_rs2; // @[RocketCore.scala 236:20]
  wire [4:0] ibuf_io_inst_0_bits_inst_rs3; // @[RocketCore.scala 236:20]
  wire [31:0] ibuf_io_inst_0_bits_raw; // @[RocketCore.scala 236:20]
  wire [29:0] ibuf_io_covSum; // @[RocketCore.scala 236:20]
  wire  ibuf_metaAssert; // @[RocketCore.scala 236:20]
  wire  ibuf_metaReset; // @[RocketCore.scala 236:20]
  reg [63:0] _T_760 [0:30]; // @[RocketCore.scala 932:23]
  reg [63:0] _RAND_0;
  wire [63:0] _T_760__T_767_data; // @[RocketCore.scala 932:23]
  wire [4:0] _T_760__T_767_addr; // @[RocketCore.scala 932:23]
  reg [63:0] _RAND_1;
  wire [63:0] _T_760__T_775_data; // @[RocketCore.scala 932:23]
  wire [4:0] _T_760__T_775_addr; // @[RocketCore.scala 932:23]
  reg [63:0] _RAND_2;
  wire [63:0] _T_760__T_1499_data; // @[RocketCore.scala 932:23]
  wire [4:0] _T_760__T_1499_addr; // @[RocketCore.scala 932:23]
  wire  _T_760__T_1499_mask; // @[RocketCore.scala 932:23]
  wire  _T_760__T_1499_en; // @[RocketCore.scala 932:23]
  wire  csr_clock; // @[RocketCore.scala 257:19]
  wire  csr_reset; // @[RocketCore.scala 257:19]
  wire  csr_io_ungated_clock; // @[RocketCore.scala 257:19]
  wire  csr_io_interrupts_debug; // @[RocketCore.scala 257:19]
  wire  csr_io_interrupts_mtip; // @[RocketCore.scala 257:19]
  wire  csr_io_interrupts_msip; // @[RocketCore.scala 257:19]
  wire  csr_io_interrupts_meip; // @[RocketCore.scala 257:19]
  wire  csr_io_interrupts_seip; // @[RocketCore.scala 257:19]
  wire [1:0] csr_io_hartid; // @[RocketCore.scala 257:19]
  wire [11:0] csr_io_rw_addr; // @[RocketCore.scala 257:19]
  wire [2:0] csr_io_rw_cmd; // @[RocketCore.scala 257:19]
  wire [63:0] csr_io_rw_rdata; // @[RocketCore.scala 257:19]
  wire [63:0] csr_io_rw_wdata; // @[RocketCore.scala 257:19]
  wire  csr_io_pcode_req_valid; // @[RocketCore.scala 257:19]
  wire [1:0] csr_io_pcode_req_bits_id; // @[RocketCore.scala 257:19]
  wire [19:0] csr_io_pcode_req_bits_value_base; // @[RocketCore.scala 257:19]
  wire [9:0] csr_io_pcode_req_bits_value_mask; // @[RocketCore.scala 257:19]
  wire  csr_io_pcode_req_bits_value_valid; // @[RocketCore.scala 257:19]
  wire  csr_io_pcode_req_bits_value_locked; // @[RocketCore.scala 257:19]
  wire [26:0] csr_io_vpoffset_req_bits_value; // @[RocketCore.scala 257:19]
  wire [11:0] csr_io_decode_0_csr; // @[RocketCore.scala 257:19]
  wire  csr_io_decode_0_fp_illegal; // @[RocketCore.scala 257:19]
  wire  csr_io_decode_0_fp_csr; // @[RocketCore.scala 257:19]
  wire  csr_io_decode_0_read_illegal; // @[RocketCore.scala 257:19]
  wire  csr_io_decode_0_write_illegal; // @[RocketCore.scala 257:19]
  wire  csr_io_decode_0_write_flush; // @[RocketCore.scala 257:19]
  wire  csr_io_decode_0_system_illegal; // @[RocketCore.scala 257:19]
  wire  csr_io_csr_stall; // @[RocketCore.scala 257:19]
  wire  csr_io_eret; // @[RocketCore.scala 257:19]
  wire  csr_io_singleStep; // @[RocketCore.scala 257:19]
  wire  csr_io_status_debug; // @[RocketCore.scala 257:19]
  wire [31:0] csr_io_status_isa; // @[RocketCore.scala 257:19]
  wire [1:0] csr_io_status_dprv; // @[RocketCore.scala 257:19]
  wire [1:0] csr_io_status_prv; // @[RocketCore.scala 257:19]
  wire  csr_io_status_sd; // @[RocketCore.scala 257:19]
  wire [26:0] csr_io_status_zero2; // @[RocketCore.scala 257:19]
  wire [1:0] csr_io_status_sxl; // @[RocketCore.scala 257:19]
  wire [1:0] csr_io_status_uxl; // @[RocketCore.scala 257:19]
  wire  csr_io_status_sd_rv32; // @[RocketCore.scala 257:19]
  wire [7:0] csr_io_status_zero1; // @[RocketCore.scala 257:19]
  wire  csr_io_status_tsr; // @[RocketCore.scala 257:19]
  wire  csr_io_status_tw; // @[RocketCore.scala 257:19]
  wire  csr_io_status_tvm; // @[RocketCore.scala 257:19]
  wire  csr_io_status_mxr; // @[RocketCore.scala 257:19]
  wire  csr_io_status_sum; // @[RocketCore.scala 257:19]
  wire  csr_io_status_mprv; // @[RocketCore.scala 257:19]
  wire [1:0] csr_io_status_xs; // @[RocketCore.scala 257:19]
  wire [1:0] csr_io_status_fs; // @[RocketCore.scala 257:19]
  wire [1:0] csr_io_status_mpp; // @[RocketCore.scala 257:19]
  wire [1:0] csr_io_status_hpp; // @[RocketCore.scala 257:19]
  wire  csr_io_status_spp; // @[RocketCore.scala 257:19]
  wire  csr_io_status_mpie; // @[RocketCore.scala 257:19]
  wire  csr_io_status_hpie; // @[RocketCore.scala 257:19]
  wire  csr_io_status_spie; // @[RocketCore.scala 257:19]
  wire  csr_io_status_upie; // @[RocketCore.scala 257:19]
  wire  csr_io_status_mie; // @[RocketCore.scala 257:19]
  wire  csr_io_status_hie; // @[RocketCore.scala 257:19]
  wire  csr_io_status_sie; // @[RocketCore.scala 257:19]
  wire  csr_io_status_uie; // @[RocketCore.scala 257:19]
  wire [3:0] csr_io_ptbr_mode; // @[RocketCore.scala 257:19]
  wire [43:0] csr_io_ptbr_ppn; // @[RocketCore.scala 257:19]
  wire [39:0] csr_io_evec; // @[RocketCore.scala 257:19]
  wire  csr_io_exception; // @[RocketCore.scala 257:19]
  wire  csr_io_retire; // @[RocketCore.scala 257:19]
  wire [63:0] csr_io_cause; // @[RocketCore.scala 257:19]
  wire [39:0] csr_io_pc; // @[RocketCore.scala 257:19]
  wire [39:0] csr_io_tval; // @[RocketCore.scala 257:19]
  wire [2:0] csr_io_fcsr_rm; // @[RocketCore.scala 257:19]
  wire  csr_io_fcsr_flags_valid; // @[RocketCore.scala 257:19]
  wire [4:0] csr_io_fcsr_flags_bits; // @[RocketCore.scala 257:19]
  wire  csr_io_interrupt; // @[RocketCore.scala 257:19]
  wire [63:0] csr_io_interrupt_cause; // @[RocketCore.scala 257:19]
  wire  csr_io_bp_0_control_action; // @[RocketCore.scala 257:19]
  wire [1:0] csr_io_bp_0_control_tmatch; // @[RocketCore.scala 257:19]
  wire  csr_io_bp_0_control_m; // @[RocketCore.scala 257:19]
  wire  csr_io_bp_0_control_s; // @[RocketCore.scala 257:19]
  wire  csr_io_bp_0_control_u; // @[RocketCore.scala 257:19]
  wire  csr_io_bp_0_control_x; // @[RocketCore.scala 257:19]
  wire  csr_io_bp_0_control_w; // @[RocketCore.scala 257:19]
  wire  csr_io_bp_0_control_r; // @[RocketCore.scala 257:19]
  wire [38:0] csr_io_bp_0_address; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_0_cfg_l; // @[RocketCore.scala 257:19]
  wire [1:0] csr_io_pmp_0_cfg_a; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_0_cfg_x; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_0_cfg_w; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_0_cfg_r; // @[RocketCore.scala 257:19]
  wire [29:0] csr_io_pmp_0_addr; // @[RocketCore.scala 257:19]
  wire [31:0] csr_io_pmp_0_mask; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_1_cfg_l; // @[RocketCore.scala 257:19]
  wire [1:0] csr_io_pmp_1_cfg_a; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_1_cfg_x; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_1_cfg_w; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_1_cfg_r; // @[RocketCore.scala 257:19]
  wire [29:0] csr_io_pmp_1_addr; // @[RocketCore.scala 257:19]
  wire [31:0] csr_io_pmp_1_mask; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_2_cfg_l; // @[RocketCore.scala 257:19]
  wire [1:0] csr_io_pmp_2_cfg_a; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_2_cfg_x; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_2_cfg_w; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_2_cfg_r; // @[RocketCore.scala 257:19]
  wire [29:0] csr_io_pmp_2_addr; // @[RocketCore.scala 257:19]
  wire [31:0] csr_io_pmp_2_mask; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_3_cfg_l; // @[RocketCore.scala 257:19]
  wire [1:0] csr_io_pmp_3_cfg_a; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_3_cfg_x; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_3_cfg_w; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_3_cfg_r; // @[RocketCore.scala 257:19]
  wire [29:0] csr_io_pmp_3_addr; // @[RocketCore.scala 257:19]
  wire [31:0] csr_io_pmp_3_mask; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_4_cfg_l; // @[RocketCore.scala 257:19]
  wire [1:0] csr_io_pmp_4_cfg_a; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_4_cfg_x; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_4_cfg_w; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_4_cfg_r; // @[RocketCore.scala 257:19]
  wire [29:0] csr_io_pmp_4_addr; // @[RocketCore.scala 257:19]
  wire [31:0] csr_io_pmp_4_mask; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_5_cfg_l; // @[RocketCore.scala 257:19]
  wire [1:0] csr_io_pmp_5_cfg_a; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_5_cfg_x; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_5_cfg_w; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_5_cfg_r; // @[RocketCore.scala 257:19]
  wire [29:0] csr_io_pmp_5_addr; // @[RocketCore.scala 257:19]
  wire [31:0] csr_io_pmp_5_mask; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_6_cfg_l; // @[RocketCore.scala 257:19]
  wire [1:0] csr_io_pmp_6_cfg_a; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_6_cfg_x; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_6_cfg_w; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_6_cfg_r; // @[RocketCore.scala 257:19]
  wire [29:0] csr_io_pmp_6_addr; // @[RocketCore.scala 257:19]
  wire [31:0] csr_io_pmp_6_mask; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_7_cfg_l; // @[RocketCore.scala 257:19]
  wire [1:0] csr_io_pmp_7_cfg_a; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_7_cfg_x; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_7_cfg_w; // @[RocketCore.scala 257:19]
  wire  csr_io_pmp_7_cfg_r; // @[RocketCore.scala 257:19]
  wire [29:0] csr_io_pmp_7_addr; // @[RocketCore.scala 257:19]
  wire [31:0] csr_io_pmp_7_mask; // @[RocketCore.scala 257:19]
  wire [29:0] csr_io_covSum; // @[RocketCore.scala 257:19]
  wire  csr_metaAssert; // @[RocketCore.scala 257:19]
  wire  csr_metaReset; // @[RocketCore.scala 257:19]
  wire  bpu_io_status_debug; // @[RocketCore.scala 302:19]
  wire [1:0] bpu_io_status_prv; // @[RocketCore.scala 302:19]
  wire  bpu_io_bp_0_control_action; // @[RocketCore.scala 302:19]
  wire [1:0] bpu_io_bp_0_control_tmatch; // @[RocketCore.scala 302:19]
  wire  bpu_io_bp_0_control_m; // @[RocketCore.scala 302:19]
  wire  bpu_io_bp_0_control_s; // @[RocketCore.scala 302:19]
  wire  bpu_io_bp_0_control_u; // @[RocketCore.scala 302:19]
  wire  bpu_io_bp_0_control_x; // @[RocketCore.scala 302:19]
  wire  bpu_io_bp_0_control_w; // @[RocketCore.scala 302:19]
  wire  bpu_io_bp_0_control_r; // @[RocketCore.scala 302:19]
  wire [38:0] bpu_io_bp_0_address; // @[RocketCore.scala 302:19]
  wire [38:0] bpu_io_pc; // @[RocketCore.scala 302:19]
  wire [38:0] bpu_io_ea; // @[RocketCore.scala 302:19]
  wire  bpu_io_xcpt_if; // @[RocketCore.scala 302:19]
  wire  bpu_io_xcpt_ld; // @[RocketCore.scala 302:19]
  wire  bpu_io_xcpt_st; // @[RocketCore.scala 302:19]
  wire  bpu_io_debug_if; // @[RocketCore.scala 302:19]
  wire  bpu_io_debug_ld; // @[RocketCore.scala 302:19]
  wire  bpu_io_debug_st; // @[RocketCore.scala 302:19]
  wire [29:0] bpu_io_covSum; // @[RocketCore.scala 302:19]
  wire  bpu_metaAssert; // @[RocketCore.scala 302:19]
  wire  alu_io_dw; // @[RocketCore.scala 361:19]
  wire [3:0] alu_io_fn; // @[RocketCore.scala 361:19]
  wire [63:0] alu_io_in2; // @[RocketCore.scala 361:19]
  wire [63:0] alu_io_in1; // @[RocketCore.scala 361:19]
  wire [63:0] alu_io_out; // @[RocketCore.scala 361:19]
  wire [63:0] alu_io_adder_out; // @[RocketCore.scala 361:19]
  wire  alu_io_cmp_out; // @[RocketCore.scala 361:19]
  wire [29:0] alu_io_covSum; // @[RocketCore.scala 361:19]
  wire  alu_metaAssert; // @[RocketCore.scala 361:19]
  wire  div_clock; // @[RocketCore.scala 376:19]
  wire  div_reset; // @[RocketCore.scala 376:19]
  wire  div_io_req_ready; // @[RocketCore.scala 376:19]
  wire  div_io_req_valid; // @[RocketCore.scala 376:19]
  wire [3:0] div_io_req_bits_fn; // @[RocketCore.scala 376:19]
  wire  div_io_req_bits_dw; // @[RocketCore.scala 376:19]
  wire [63:0] div_io_req_bits_in1; // @[RocketCore.scala 376:19]
  wire [63:0] div_io_req_bits_in2; // @[RocketCore.scala 376:19]
  wire [4:0] div_io_req_bits_tag; // @[RocketCore.scala 376:19]
  wire  div_io_kill; // @[RocketCore.scala 376:19]
  wire  div_io_resp_ready; // @[RocketCore.scala 376:19]
  wire  div_io_resp_valid; // @[RocketCore.scala 376:19]
  wire [63:0] div_io_resp_bits_data; // @[RocketCore.scala 376:19]
  wire [4:0] div_io_resp_bits_tag; // @[RocketCore.scala 376:19]
  wire [29:0] div_io_covSum; // @[RocketCore.scala 376:19]
  wire  div_metaAssert; // @[RocketCore.scala 376:19]
  wire  div_metaReset; // @[RocketCore.scala 376:19]
  reg  imem_might_request_reg; // @[RocketCore.scala 112:35]
  reg [31:0] _RAND_3;
  reg  ex_ctrl_fp; // @[RocketCore.scala 182:20]
  reg [31:0] _RAND_4;
  reg  ex_ctrl_branch; // @[RocketCore.scala 182:20]
  reg [31:0] _RAND_5;
  reg  ex_ctrl_jal; // @[RocketCore.scala 182:20]
  reg [31:0] _RAND_6;
  reg  ex_ctrl_jalr; // @[RocketCore.scala 182:20]
  reg [31:0] _RAND_7;
  reg  ex_ctrl_rxs2; // @[RocketCore.scala 182:20]
  reg [31:0] _RAND_8;
  reg [1:0] ex_ctrl_sel_alu2; // @[RocketCore.scala 182:20]
  reg [31:0] _RAND_9;
  reg [1:0] ex_ctrl_sel_alu1; // @[RocketCore.scala 182:20]
  reg [31:0] _RAND_10;
  reg [2:0] ex_ctrl_sel_imm; // @[RocketCore.scala 182:20]
  reg [31:0] _RAND_11;
  reg  ex_ctrl_alu_dw; // @[RocketCore.scala 182:20]
  reg [31:0] _RAND_12;
  reg [3:0] ex_ctrl_alu_fn; // @[RocketCore.scala 182:20]
  reg [31:0] _RAND_13;
  reg  ex_ctrl_mem; // @[RocketCore.scala 182:20]
  reg [31:0] _RAND_14;
  reg [4:0] ex_ctrl_mem_cmd; // @[RocketCore.scala 182:20]
  reg [31:0] _RAND_15;
  reg [2:0] ex_ctrl_mem_type; // @[RocketCore.scala 182:20]
  reg [31:0] _RAND_16;
  reg  ex_ctrl_wfd; // @[RocketCore.scala 182:20]
  reg [31:0] _RAND_17;
  reg  ex_ctrl_div; // @[RocketCore.scala 182:20]
  reg [31:0] _RAND_18;
  reg  ex_ctrl_wxd; // @[RocketCore.scala 182:20]
  reg [31:0] _RAND_19;
  reg [2:0] ex_ctrl_csr; // @[RocketCore.scala 182:20]
  reg [31:0] _RAND_20;
  reg  ex_ctrl_fence_i; // @[RocketCore.scala 182:20]
  reg [31:0] _RAND_21;
  reg  mem_ctrl_fp; // @[RocketCore.scala 183:21]
  reg [31:0] _RAND_22;
  reg  mem_ctrl_branch; // @[RocketCore.scala 183:21]
  reg [31:0] _RAND_23;
  reg  mem_ctrl_jal; // @[RocketCore.scala 183:21]
  reg [31:0] _RAND_24;
  reg  mem_ctrl_jalr; // @[RocketCore.scala 183:21]
  reg [31:0] _RAND_25;
  reg  mem_ctrl_mem; // @[RocketCore.scala 183:21]
  reg [31:0] _RAND_26;
  reg [2:0] mem_ctrl_mem_type; // @[RocketCore.scala 183:21]
  reg [31:0] _RAND_27;
  reg  mem_ctrl_wfd; // @[RocketCore.scala 183:21]
  reg [31:0] _RAND_28;
  reg  mem_ctrl_div; // @[RocketCore.scala 183:21]
  reg [31:0] _RAND_29;
  reg  mem_ctrl_wxd; // @[RocketCore.scala 183:21]
  reg [31:0] _RAND_30;
  reg [2:0] mem_ctrl_csr; // @[RocketCore.scala 183:21]
  reg [31:0] _RAND_31;
  reg  mem_ctrl_fence_i; // @[RocketCore.scala 183:21]
  reg [31:0] _RAND_32;
  reg  wb_ctrl_mem; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_33;
  reg [2:0] wb_ctrl_mem_type; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_34;
  reg  wb_ctrl_wfd; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_35;
  reg  wb_ctrl_div; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_36;
  reg  wb_ctrl_wxd; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_37;
  reg [2:0] wb_ctrl_csr; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_38;
  reg  wb_ctrl_fence_i; // @[RocketCore.scala 184:20]
  reg [31:0] _RAND_39;
  reg  ex_reg_xcpt_interrupt; // @[RocketCore.scala 186:35]
  reg [31:0] _RAND_40;
  reg  ex_reg_valid; // @[RocketCore.scala 187:35]
  reg [31:0] _RAND_41;
  reg  ex_reg_rvc; // @[RocketCore.scala 188:35]
  reg [31:0] _RAND_42;
  reg [4:0] ex_reg_btb_resp_entry; // @[RocketCore.scala 189:35]
  reg [31:0] _RAND_43;
  reg [7:0] ex_reg_btb_resp_bht_history; // @[RocketCore.scala 189:35]
  reg [31:0] _RAND_44;
  reg  ex_reg_xcpt; // @[RocketCore.scala 190:35]
  reg [31:0] _RAND_45;
  reg  ex_reg_flush_pipe; // @[RocketCore.scala 191:35]
  reg [31:0] _RAND_46;
  reg  ex_reg_load_use; // @[RocketCore.scala 192:35]
  reg [31:0] _RAND_47;
  reg [63:0] ex_reg_cause; // @[RocketCore.scala 193:35]
  reg [63:0] _RAND_48;
  reg  ex_reg_replay; // @[RocketCore.scala 194:26]
  reg [31:0] _RAND_49;
  reg [39:0] ex_reg_pc; // @[RocketCore.scala 195:22]
  reg [63:0] _RAND_50;
  reg [31:0] ex_reg_inst; // @[RocketCore.scala 196:24]
  reg [31:0] _RAND_51;
  reg  mem_reg_xcpt_interrupt; // @[RocketCore.scala 199:36]
  reg [31:0] _RAND_52;
  reg  mem_reg_valid; // @[RocketCore.scala 200:36]
  reg [31:0] _RAND_53;
  reg  mem_reg_rvc; // @[RocketCore.scala 201:36]
  reg [31:0] _RAND_54;
  reg [4:0] mem_reg_btb_resp_entry; // @[RocketCore.scala 202:36]
  reg [31:0] _RAND_55;
  reg [7:0] mem_reg_btb_resp_bht_history; // @[RocketCore.scala 202:36]
  reg [31:0] _RAND_56;
  reg  mem_reg_xcpt; // @[RocketCore.scala 203:36]
  reg [31:0] _RAND_57;
  reg  mem_reg_replay; // @[RocketCore.scala 204:36]
  reg [31:0] _RAND_58;
  reg  mem_reg_flush_pipe; // @[RocketCore.scala 205:36]
  reg [31:0] _RAND_59;
  reg [63:0] mem_reg_cause; // @[RocketCore.scala 206:36]
  reg [63:0] _RAND_60;
  reg  mem_reg_slow_bypass; // @[RocketCore.scala 207:36]
  reg [31:0] _RAND_61;
  reg  mem_reg_load; // @[RocketCore.scala 208:36]
  reg [31:0] _RAND_62;
  reg  mem_reg_store; // @[RocketCore.scala 209:36]
  reg [31:0] _RAND_63;
  reg  mem_reg_sfence; // @[RocketCore.scala 210:27]
  reg [31:0] _RAND_64;
  reg [39:0] mem_reg_pc; // @[RocketCore.scala 211:23]
  reg [63:0] _RAND_65;
  reg [31:0] mem_reg_inst; // @[RocketCore.scala 212:25]
  reg [31:0] _RAND_66;
  reg [63:0] mem_reg_wdata; // @[RocketCore.scala 214:26]
  reg [63:0] _RAND_67;
  reg [63:0] mem_reg_rs2; // @[RocketCore.scala 215:24]
  reg [63:0] _RAND_68;
  reg  mem_br_taken; // @[RocketCore.scala 216:25]
  reg [31:0] _RAND_69;
  reg  wb_reg_valid; // @[RocketCore.scala 219:35]
  reg [31:0] _RAND_70;
  reg  wb_reg_xcpt; // @[RocketCore.scala 220:35]
  reg [31:0] _RAND_71;
  reg  wb_reg_replay; // @[RocketCore.scala 221:35]
  reg [31:0] _RAND_72;
  reg  wb_reg_flush_pipe; // @[RocketCore.scala 222:35]
  reg [31:0] _RAND_73;
  reg [63:0] wb_reg_cause; // @[RocketCore.scala 223:35]
  reg [63:0] _RAND_74;
  reg  wb_reg_sfence; // @[RocketCore.scala 224:26]
  reg [31:0] _RAND_75;
  reg [39:0] wb_reg_pc; // @[RocketCore.scala 225:22]
  reg [63:0] _RAND_76;
  reg [31:0] wb_reg_inst; // @[RocketCore.scala 226:24]
  reg [31:0] _RAND_77;
  reg [63:0] wb_reg_wdata; // @[RocketCore.scala 228:25]
  reg [63:0] _RAND_78;
  wire  replay_wb_common; // @[RocketCore.scala 585:42]
  wire  _T_1437; // @[RocketCore.scala 564:19]
  wire  _T_1438; // @[RocketCore.scala 564:34]
  wire  _T_1449; // @[RocketCore.scala 892:26]
  wire  _T_1440; // @[RocketCore.scala 565:34]
  wire  _T_1450; // @[RocketCore.scala 892:26]
  wire  _T_1442; // @[RocketCore.scala 566:34]
  wire  _T_1451; // @[RocketCore.scala 892:26]
  wire  _T_1444; // @[RocketCore.scala 567:34]
  wire  _T_1452; // @[RocketCore.scala 892:26]
  wire  _T_1446; // @[RocketCore.scala 568:34]
  wire  _T_1453; // @[RocketCore.scala 892:26]
  wire  _T_1448; // @[RocketCore.scala 569:34]
  wire  wb_xcpt; // @[RocketCore.scala 892:26]
  wire  _T_1475; // @[RocketCore.scala 588:27]
  wire  _T_1476; // @[RocketCore.scala 588:38]
  wire  take_pc_wb; // @[RocketCore.scala 588:53]
  wire  _T_1109; // @[RocketCore.scala 447:34]
  wire  ex_pc_valid; // @[RocketCore.scala 447:51]
  wire  _T_1282; // @[RocketCore.scala 470:36]
  wire [24:0] a; // @[RocketCore.scala 906:23]
  wire  _T_1284; // @[RocketCore.scala 907:21]
  wire  _T_1285; // @[RocketCore.scala 907:34]
  wire  _T_1286; // @[RocketCore.scala 907:29]
  wire  msb; // @[RocketCore.scala 907:18]
  wire [39:0] _T_1292; // @[RocketCore.scala 470:106]
  wire  _T_1152; // @[RocketCore.scala 467:25]
  wire  _T_1155; // @[RocketCore.scala 954:53]
  wire  _T_1210; // @[Cat.scala 30:58]
  wire [10:0] _T_1209; // @[Cat.scala 30:58]
  wire [7:0] _T_1207; // @[Cat.scala 30:58]
  wire  _T_1206; // @[Cat.scala 30:58]
  wire [31:0] _T_1214; // @[RocketCore.scala 968:53]
  wire [7:0] _T_1269; // @[Cat.scala 30:58]
  wire  _T_1268; // @[Cat.scala 30:58]
  wire [31:0] _T_1276; // @[RocketCore.scala 968:53]
  wire [3:0] _T_1277; // @[RocketCore.scala 469:8]
  wire [31:0] _T_1278; // @[RocketCore.scala 468:8]
  wire [31:0] _T_1279; // @[RocketCore.scala 467:8]
  wire [39:0] _GEN_235; // @[RocketCore.scala 466:41]
  wire [39:0] mem_br_target; // @[RocketCore.scala 466:41]
  wire [39:0] _T_1293; // @[RocketCore.scala 470:21]
  wire [39:0] mem_npc; // @[RocketCore.scala 470:141]
  wire  _T_1296; // @[RocketCore.scala 472:30]
  wire  _T_1297; // @[RocketCore.scala 473:31]
  wire  _T_1298; // @[RocketCore.scala 473:62]
  wire  _T_1299; // @[RocketCore.scala 473:8]
  wire  mem_wrong_npc; // @[RocketCore.scala 472:8]
  wire  _T_1315; // @[RocketCore.scala 480:54]
  wire  take_pc_mem; // @[RocketCore.scala 480:32]
  wire  take_pc_mem_wb; // @[RocketCore.scala 232:35]
  wire [31:0] _T_309; // @[Decode.scala 14:65]
  wire  _T_310; // @[Decode.scala 14:121]
  wire [31:0] _T_311; // @[Decode.scala 14:65]
  wire  _T_312; // @[Decode.scala 14:121]
  wire [31:0] _T_313; // @[Decode.scala 14:65]
  wire  _T_314; // @[Decode.scala 14:121]
  wire [31:0] _T_315; // @[Decode.scala 14:65]
  wire  _T_316; // @[Decode.scala 14:121]
  wire [31:0] _T_317; // @[Decode.scala 14:65]
  wire  _T_318; // @[Decode.scala 14:121]
  wire [31:0] _T_319; // @[Decode.scala 14:65]
  wire  _T_320; // @[Decode.scala 14:121]
  wire [31:0] _T_321; // @[Decode.scala 14:65]
  wire  _T_322; // @[Decode.scala 14:121]
  wire [31:0] _T_323; // @[Decode.scala 14:65]
  wire  _T_324; // @[Decode.scala 14:121]
  wire [31:0] _T_325; // @[Decode.scala 14:65]
  wire  _T_326; // @[Decode.scala 14:121]
  wire [31:0] _T_327; // @[Decode.scala 14:65]
  wire  _T_328; // @[Decode.scala 14:121]
  wire [31:0] _T_329; // @[Decode.scala 14:65]
  wire  _T_330; // @[Decode.scala 14:121]
  wire [31:0] _T_331; // @[Decode.scala 14:65]
  wire  _T_332; // @[Decode.scala 14:121]
  wire [31:0] _T_333; // @[Decode.scala 14:65]
  wire  _T_334; // @[Decode.scala 14:121]
  wire [31:0] _T_335; // @[Decode.scala 14:65]
  wire  _T_336; // @[Decode.scala 14:121]
  wire [31:0] _T_337; // @[Decode.scala 14:65]
  wire  _T_338; // @[Decode.scala 14:121]
  wire  _T_340; // @[Decode.scala 14:121]
  wire [31:0] _T_341; // @[Decode.scala 14:65]
  wire  _T_342; // @[Decode.scala 14:121]
  wire  _T_344; // @[Decode.scala 14:121]
  wire [31:0] _T_345; // @[Decode.scala 14:65]
  wire  _T_346; // @[Decode.scala 14:121]
  wire [31:0] _T_347; // @[Decode.scala 14:65]
  wire  _T_348; // @[Decode.scala 14:121]
  wire  _T_350; // @[Decode.scala 14:121]
  wire [31:0] _T_351; // @[Decode.scala 14:65]
  wire  _T_352; // @[Decode.scala 14:121]
  wire [31:0] _T_353; // @[Decode.scala 14:65]
  wire  _T_354; // @[Decode.scala 14:121]
  wire [31:0] _T_355; // @[Decode.scala 14:65]
  wire  _T_356; // @[Decode.scala 14:121]
  wire [31:0] _T_357; // @[Decode.scala 14:65]
  wire  _T_358; // @[Decode.scala 14:121]
  wire  _T_359; // @[Decode.scala 14:121]
  wire [31:0] _T_360; // @[Decode.scala 14:65]
  wire  _T_361; // @[Decode.scala 14:121]
  wire [31:0] _T_362; // @[Decode.scala 14:65]
  wire  _T_363; // @[Decode.scala 14:121]
  wire [31:0] _T_364; // @[Decode.scala 14:65]
  wire  _T_365; // @[Decode.scala 14:121]
  wire [31:0] _T_366; // @[Decode.scala 14:65]
  wire  _T_367; // @[Decode.scala 14:121]
  wire [31:0] _T_368; // @[Decode.scala 14:65]
  wire  _T_369; // @[Decode.scala 14:121]
  wire  _T_371; // @[Decode.scala 14:121]
  wire [31:0] _T_372; // @[Decode.scala 14:65]
  wire  _T_373; // @[Decode.scala 14:121]
  wire  _T_374; // @[Decode.scala 14:121]
  wire [31:0] _T_375; // @[Decode.scala 14:65]
  wire  _T_376; // @[Decode.scala 14:121]
  wire [31:0] _T_377; // @[Decode.scala 14:65]
  wire  _T_378; // @[Decode.scala 14:121]
  wire [31:0] _T_379; // @[Decode.scala 14:65]
  wire  _T_380; // @[Decode.scala 14:121]
  wire [31:0] _T_381; // @[Decode.scala 14:65]
  wire  _T_382; // @[Decode.scala 14:121]
  wire [31:0] _T_383; // @[Decode.scala 14:65]
  wire  _T_384; // @[Decode.scala 14:121]
  wire [31:0] _T_385; // @[Decode.scala 14:65]
  wire  _T_386; // @[Decode.scala 14:121]
  wire [31:0] _T_387; // @[Decode.scala 14:65]
  wire  _T_388; // @[Decode.scala 14:121]
  wire  _T_390; // @[Decode.scala 15:30]
  wire  _T_391; // @[Decode.scala 15:30]
  wire  _T_392; // @[Decode.scala 15:30]
  wire  _T_393; // @[Decode.scala 15:30]
  wire  _T_394; // @[Decode.scala 15:30]
  wire  _T_395; // @[Decode.scala 15:30]
  wire  _T_396; // @[Decode.scala 15:30]
  wire  _T_397; // @[Decode.scala 15:30]
  wire  _T_398; // @[Decode.scala 15:30]
  wire  _T_399; // @[Decode.scala 15:30]
  wire  _T_400; // @[Decode.scala 15:30]
  wire  _T_401; // @[Decode.scala 15:30]
  wire  _T_402; // @[Decode.scala 15:30]
  wire  _T_403; // @[Decode.scala 15:30]
  wire  _T_404; // @[Decode.scala 15:30]
  wire  _T_405; // @[Decode.scala 15:30]
  wire  _T_406; // @[Decode.scala 15:30]
  wire  _T_407; // @[Decode.scala 15:30]
  wire  _T_408; // @[Decode.scala 15:30]
  wire  _T_409; // @[Decode.scala 15:30]
  wire  _T_410; // @[Decode.scala 15:30]
  wire  _T_411; // @[Decode.scala 15:30]
  wire  _T_412; // @[Decode.scala 15:30]
  wire  _T_413; // @[Decode.scala 15:30]
  wire  _T_414; // @[Decode.scala 15:30]
  wire  _T_415; // @[Decode.scala 15:30]
  wire  _T_416; // @[Decode.scala 15:30]
  wire  _T_417; // @[Decode.scala 15:30]
  wire  _T_418; // @[Decode.scala 15:30]
  wire  _T_419; // @[Decode.scala 15:30]
  wire  _T_420; // @[Decode.scala 15:30]
  wire  _T_421; // @[Decode.scala 15:30]
  wire  _T_422; // @[Decode.scala 15:30]
  wire  _T_423; // @[Decode.scala 15:30]
  wire  _T_424; // @[Decode.scala 15:30]
  wire  _T_425; // @[Decode.scala 15:30]
  wire  _T_426; // @[Decode.scala 15:30]
  wire  _T_427; // @[Decode.scala 15:30]
  wire  _T_428; // @[Decode.scala 15:30]
  wire  id_ctrl_legal; // @[Decode.scala 15:30]
  wire [31:0] _T_430; // @[Decode.scala 14:65]
  wire  _T_431; // @[Decode.scala 14:121]
  wire [31:0] _T_432; // @[Decode.scala 14:65]
  wire  _T_433; // @[Decode.scala 14:121]
  wire  id_ctrl_fp; // @[Decode.scala 15:30]
  wire [31:0] _T_436; // @[Decode.scala 14:65]
  wire  id_ctrl_branch; // @[Decode.scala 14:121]
  wire [31:0] _T_439; // @[Decode.scala 14:65]
  wire  id_ctrl_jal; // @[Decode.scala 14:121]
  wire [31:0] _T_442; // @[Decode.scala 14:65]
  wire  id_ctrl_jalr; // @[Decode.scala 14:121]
  wire [31:0] _T_445; // @[Decode.scala 14:65]
  wire  _T_446; // @[Decode.scala 14:121]
  wire [31:0] _T_447; // @[Decode.scala 14:65]
  wire  _T_448; // @[Decode.scala 14:121]
  wire [31:0] _T_449; // @[Decode.scala 14:65]
  wire  _T_450; // @[Decode.scala 14:121]
  wire [31:0] _T_451; // @[Decode.scala 14:65]
  wire  _T_452; // @[Decode.scala 14:121]
  wire  _T_454; // @[Decode.scala 15:30]
  wire  _T_455; // @[Decode.scala 15:30]
  wire  id_ctrl_rxs2; // @[Decode.scala 15:30]
  wire [31:0] _T_457; // @[Decode.scala 14:65]
  wire  _T_458; // @[Decode.scala 14:121]
  wire [31:0] _T_459; // @[Decode.scala 14:65]
  wire  _T_460; // @[Decode.scala 14:121]
  wire [31:0] _T_461; // @[Decode.scala 14:65]
  wire  _T_462; // @[Decode.scala 14:121]
  wire [31:0] _T_463; // @[Decode.scala 14:65]
  wire  _T_464; // @[Decode.scala 14:121]
  wire [31:0] _T_465; // @[Decode.scala 14:65]
  wire  _T_466; // @[Decode.scala 14:121]
  wire  _T_468; // @[Decode.scala 15:30]
  wire  _T_469; // @[Decode.scala 15:30]
  wire  _T_470; // @[Decode.scala 15:30]
  wire  id_ctrl_rxs1; // @[Decode.scala 15:30]
  wire [31:0] _T_472; // @[Decode.scala 14:65]
  wire  _T_473; // @[Decode.scala 14:121]
  wire [31:0] _T_474; // @[Decode.scala 14:65]
  wire  _T_475; // @[Decode.scala 14:121]
  wire [31:0] _T_476; // @[Decode.scala 14:65]
  wire  _T_477; // @[Decode.scala 14:121]
  wire [31:0] _T_478; // @[Decode.scala 14:65]
  wire  _T_479; // @[Decode.scala 14:121]
  wire [31:0] _T_480; // @[Decode.scala 14:65]
  wire  _T_481; // @[Decode.scala 14:121]
  wire  _T_483; // @[Decode.scala 15:30]
  wire  _T_484; // @[Decode.scala 15:30]
  wire  _T_485; // @[Decode.scala 15:30]
  wire  _T_486; // @[Decode.scala 15:30]
  wire  _T_488; // @[Decode.scala 14:121]
  wire [31:0] _T_489; // @[Decode.scala 14:65]
  wire  _T_490; // @[Decode.scala 14:121]
  wire [31:0] _T_491; // @[Decode.scala 14:65]
  wire  _T_492; // @[Decode.scala 14:121]
  wire  _T_494; // @[Decode.scala 15:30]
  wire  _T_495; // @[Decode.scala 15:30]
  wire  _T_496; // @[Decode.scala 15:30]
  wire [1:0] id_ctrl_sel_alu2; // @[Cat.scala 30:58]
  wire [31:0] _T_498; // @[Decode.scala 14:65]
  wire  _T_499; // @[Decode.scala 14:121]
  wire [31:0] _T_500; // @[Decode.scala 14:65]
  wire  _T_501; // @[Decode.scala 14:121]
  wire [31:0] _T_502; // @[Decode.scala 14:65]
  wire  _T_503; // @[Decode.scala 14:121]
  wire  _T_505; // @[Decode.scala 15:30]
  wire  _T_506; // @[Decode.scala 15:30]
  wire  _T_507; // @[Decode.scala 15:30]
  wire  _T_508; // @[Decode.scala 15:30]
  wire  _T_510; // @[Decode.scala 14:121]
  wire  _T_512; // @[Decode.scala 15:30]
  wire [1:0] id_ctrl_sel_alu1; // @[Cat.scala 30:58]
  wire  _T_515; // @[Decode.scala 14:121]
  wire  _T_517; // @[Decode.scala 14:121]
  wire  _T_519; // @[Decode.scala 15:30]
  wire [31:0] _T_520; // @[Decode.scala 14:65]
  wire  _T_521; // @[Decode.scala 14:121]
  wire  _T_523; // @[Decode.scala 15:30]
  wire [31:0] _T_524; // @[Decode.scala 14:65]
  wire  _T_525; // @[Decode.scala 14:121]
  wire [31:0] _T_526; // @[Decode.scala 14:65]
  wire  _T_527; // @[Decode.scala 14:121]
  wire  _T_529; // @[Decode.scala 14:121]
  wire  _T_531; // @[Decode.scala 15:30]
  wire  _T_532; // @[Decode.scala 15:30]
  wire [2:0] id_ctrl_sel_imm; // @[Cat.scala 30:58]
  wire [31:0] _T_535; // @[Decode.scala 14:65]
  wire  _T_536; // @[Decode.scala 14:121]
  wire [31:0] _T_537; // @[Decode.scala 14:65]
  wire  _T_538; // @[Decode.scala 14:121]
  wire  id_ctrl_alu_dw; // @[Decode.scala 15:30]
  wire [31:0] _T_541; // @[Decode.scala 14:65]
  wire  _T_542; // @[Decode.scala 14:121]
  wire [31:0] _T_543; // @[Decode.scala 14:65]
  wire  _T_544; // @[Decode.scala 14:121]
  wire [31:0] _T_545; // @[Decode.scala 14:65]
  wire  _T_546; // @[Decode.scala 14:121]
  wire [31:0] _T_547; // @[Decode.scala 14:65]
  wire  _T_548; // @[Decode.scala 14:121]
  wire  _T_550; // @[Decode.scala 15:30]
  wire  _T_551; // @[Decode.scala 15:30]
  wire  _T_552; // @[Decode.scala 15:30]
  wire [31:0] _T_553; // @[Decode.scala 14:65]
  wire  _T_554; // @[Decode.scala 14:121]
  wire [31:0] _T_555; // @[Decode.scala 14:65]
  wire  _T_556; // @[Decode.scala 14:121]
  wire  _T_558; // @[Decode.scala 14:121]
  wire [31:0] _T_559; // @[Decode.scala 14:65]
  wire  _T_560; // @[Decode.scala 14:121]
  wire [31:0] _T_561; // @[Decode.scala 14:65]
  wire  _T_562; // @[Decode.scala 14:121]
  wire [31:0] _T_563; // @[Decode.scala 14:65]
  wire  _T_564; // @[Decode.scala 14:121]
  wire [31:0] _T_565; // @[Decode.scala 14:65]
  wire  _T_566; // @[Decode.scala 14:121]
  wire  _T_568; // @[Decode.scala 15:30]
  wire  _T_569; // @[Decode.scala 15:30]
  wire  _T_570; // @[Decode.scala 15:30]
  wire  _T_571; // @[Decode.scala 15:30]
  wire  _T_572; // @[Decode.scala 15:30]
  wire  _T_573; // @[Decode.scala 15:30]
  wire [31:0] _T_574; // @[Decode.scala 14:65]
  wire  _T_575; // @[Decode.scala 14:121]
  wire [31:0] _T_576; // @[Decode.scala 14:65]
  wire  _T_577; // @[Decode.scala 14:121]
  wire [31:0] _T_578; // @[Decode.scala 14:65]
  wire  _T_579; // @[Decode.scala 14:121]
  wire [31:0] _T_580; // @[Decode.scala 14:65]
  wire  _T_581; // @[Decode.scala 14:121]
  wire [31:0] _T_582; // @[Decode.scala 14:65]
  wire  _T_583; // @[Decode.scala 14:121]
  wire  _T_585; // @[Decode.scala 15:30]
  wire  _T_586; // @[Decode.scala 15:30]
  wire  _T_587; // @[Decode.scala 15:30]
  wire  _T_588; // @[Decode.scala 15:30]
  wire [31:0] _T_589; // @[Decode.scala 14:65]
  wire  _T_590; // @[Decode.scala 14:121]
  wire [31:0] _T_591; // @[Decode.scala 14:65]
  wire  _T_592; // @[Decode.scala 14:121]
  wire [31:0] _T_593; // @[Decode.scala 14:65]
  wire  _T_594; // @[Decode.scala 14:121]
  wire  _T_596; // @[Decode.scala 15:30]
  wire  _T_597; // @[Decode.scala 15:30]
  wire  _T_598; // @[Decode.scala 15:30]
  wire  _T_599; // @[Decode.scala 15:30]
  wire [3:0] id_ctrl_alu_fn; // @[Cat.scala 30:58]
  wire [31:0] _T_603; // @[Decode.scala 14:65]
  wire  _T_604; // @[Decode.scala 14:121]
  wire [31:0] _T_605; // @[Decode.scala 14:65]
  wire  _T_606; // @[Decode.scala 14:121]
  wire  _T_608; // @[Decode.scala 15:30]
  wire  _T_609; // @[Decode.scala 15:30]
  wire  _T_610; // @[Decode.scala 15:30]
  wire  _T_611; // @[Decode.scala 15:30]
  wire  _T_612; // @[Decode.scala 15:30]
  wire  _T_613; // @[Decode.scala 15:30]
  wire  _T_614; // @[Decode.scala 15:30]
  wire  id_ctrl_mem; // @[Decode.scala 15:30]
  wire [31:0] _T_616; // @[Decode.scala 14:65]
  wire  _T_617; // @[Decode.scala 14:121]
  wire  _T_619; // @[Decode.scala 14:121]
  wire [31:0] _T_620; // @[Decode.scala 14:65]
  wire  _T_621; // @[Decode.scala 14:121]
  wire [31:0] _T_622; // @[Decode.scala 14:65]
  wire  _T_623; // @[Decode.scala 14:121]
  wire  _T_625; // @[Decode.scala 15:30]
  wire  _T_626; // @[Decode.scala 15:30]
  wire  _T_627; // @[Decode.scala 15:30]
  wire [31:0] _T_628; // @[Decode.scala 14:65]
  wire  _T_629; // @[Decode.scala 14:121]
  wire [31:0] _T_630; // @[Decode.scala 14:65]
  wire  _T_631; // @[Decode.scala 14:121]
  wire  _T_633; // @[Decode.scala 15:30]
  wire [31:0] _T_634; // @[Decode.scala 14:65]
  wire  _T_635; // @[Decode.scala 14:121]
  wire [31:0] _T_636; // @[Decode.scala 14:65]
  wire  _T_637; // @[Decode.scala 14:121]
  wire [31:0] _T_638; // @[Decode.scala 14:65]
  wire  _T_639; // @[Decode.scala 14:121]
  wire [31:0] _T_640; // @[Decode.scala 14:65]
  wire  _T_641; // @[Decode.scala 14:121]
  wire  _T_643; // @[Decode.scala 15:30]
  wire  _T_644; // @[Decode.scala 15:30]
  wire  _T_645; // @[Decode.scala 15:30]
  wire  _T_646; // @[Decode.scala 15:30]
  wire [31:0] _T_647; // @[Decode.scala 14:65]
  wire  _T_648; // @[Decode.scala 14:121]
  wire [4:0] id_ctrl_mem_cmd; // @[Cat.scala 30:58]
  wire [31:0] _T_655; // @[Decode.scala 14:65]
  wire  _T_656; // @[Decode.scala 14:121]
  wire [31:0] _T_658; // @[Decode.scala 14:65]
  wire  _T_659; // @[Decode.scala 14:121]
  wire  _T_661; // @[Decode.scala 15:30]
  wire [31:0] _T_662; // @[Decode.scala 14:65]
  wire  _T_663; // @[Decode.scala 14:121]
  wire [2:0] id_ctrl_mem_type; // @[Cat.scala 30:58]
  wire [31:0] _T_667; // @[Decode.scala 14:65]
  wire  _T_668; // @[Decode.scala 14:121]
  wire [31:0] _T_669; // @[Decode.scala 14:65]
  wire [31:0] _T_671; // @[Decode.scala 14:65]
  wire  id_ctrl_rfs3; // @[Decode.scala 14:121]
  wire [31:0] _T_687; // @[Decode.scala 14:65]
  wire  _T_688; // @[Decode.scala 14:121]
  wire  _T_690; // @[Decode.scala 14:121]
  wire  _T_692; // @[Decode.scala 15:30]
  wire  _T_693; // @[Decode.scala 15:30]
  wire  id_ctrl_wfd; // @[Decode.scala 15:30]
  wire [31:0] _T_695; // @[Decode.scala 14:65]
  wire  id_ctrl_div; // @[Decode.scala 14:121]
  wire  _T_699; // @[Decode.scala 14:121]
  wire  _T_701; // @[Decode.scala 14:121]
  wire [31:0] _T_702; // @[Decode.scala 14:65]
  wire  _T_703; // @[Decode.scala 14:121]
  wire [31:0] _T_704; // @[Decode.scala 14:65]
  wire  _T_705; // @[Decode.scala 14:121]
  wire [31:0] _T_706; // @[Decode.scala 14:65]
  wire  _T_707; // @[Decode.scala 14:121]
  wire [31:0] _T_708; // @[Decode.scala 14:65]
  wire  _T_709; // @[Decode.scala 14:121]
  wire [31:0] _T_710; // @[Decode.scala 14:65]
  wire  _T_711; // @[Decode.scala 14:121]
  wire  _T_713; // @[Decode.scala 15:30]
  wire  _T_714; // @[Decode.scala 15:30]
  wire  _T_715; // @[Decode.scala 15:30]
  wire  _T_716; // @[Decode.scala 15:30]
  wire  _T_717; // @[Decode.scala 15:30]
  wire  id_ctrl_wxd; // @[Decode.scala 15:30]
  wire [31:0] _T_719; // @[Decode.scala 14:65]
  wire  _T_720; // @[Decode.scala 14:121]
  wire [31:0] _T_722; // @[Decode.scala 14:65]
  wire  _T_723; // @[Decode.scala 14:121]
  wire [31:0] _T_725; // @[Decode.scala 14:65]
  wire  _T_726; // @[Decode.scala 14:121]
  wire [31:0] _T_727; // @[Decode.scala 14:65]
  wire  _T_728; // @[Decode.scala 14:121]
  wire [31:0] _T_729; // @[Decode.scala 14:65]
  wire  _T_730; // @[Decode.scala 14:121]
  wire  _T_732; // @[Decode.scala 15:30]
  wire  _T_733; // @[Decode.scala 15:30]
  wire  _T_734; // @[Decode.scala 15:30]
  wire  _T_735; // @[Decode.scala 15:30]
  wire [2:0] id_ctrl_csr; // @[Cat.scala 30:58]
  wire [31:0] _T_738; // @[Decode.scala 14:65]
  wire  id_ctrl_fence_i; // @[Decode.scala 14:121]
  wire  id_ctrl_fence; // @[Decode.scala 14:121]
  wire [31:0] _T_744; // @[Decode.scala 14:65]
  wire  id_ctrl_amo; // @[Decode.scala 14:121]
  wire [31:0] _T_747; // @[Decode.scala 14:65]
  wire  _T_748; // @[Decode.scala 14:121]
  wire [31:0] _T_749; // @[Decode.scala 14:65]
  wire  _T_750; // @[Decode.scala 14:121]
  wire [31:0] _T_751; // @[Decode.scala 14:65]
  wire  _T_752; // @[Decode.scala 14:121]
  wire  _T_754; // @[Decode.scala 15:30]
  wire  id_ctrl_dp; // @[Decode.scala 15:30]
  reg  id_reg_fence; // @[RocketCore.scala 250:25]
  reg [31:0] _RAND_79;
  wire  _T_763; // @[RocketCore.scala 939:45]
  wire [4:0] _T_765; // @[RocketCore.scala 933:44]
  wire [63:0] _T_768; // @[RocketCore.scala 939:25]
  wire [4:0] _T_773; // @[RocketCore.scala 933:44]
  wire [63:0] _T_776; // @[RocketCore.scala 939:25]
  wire  _T_847; // @[package.scala 14:47]
  wire  _T_848; // @[package.scala 14:47]
  wire  _T_849; // @[package.scala 14:47]
  wire  _T_850; // @[package.scala 14:62]
  wire  id_csr_en; // @[package.scala 14:62]
  wire  id_system_insn; // @[RocketCore.scala 259:36]
  wire  id_csr_ren; // @[RocketCore.scala 260:54]
  wire  _T_855; // @[RocketCore.scala 262:50]
  wire  id_sfence; // @[RocketCore.scala 262:31]
  wire  _T_856; // @[RocketCore.scala 263:32]
  wire  _T_858; // @[RocketCore.scala 263:64]
  wire  _T_859; // @[RocketCore.scala 263:79]
  wire  id_csr_flush; // @[RocketCore.scala 263:50]
  wire  _T_864; // @[RocketCore.scala 281:34]
  wire  _T_865; // @[RocketCore.scala 280:40]
  wire  _T_868; // @[RocketCore.scala 282:17]
  wire  _T_869; // @[RocketCore.scala 281:65]
  wire  _T_870; // @[RocketCore.scala 283:48]
  wire  _T_871; // @[RocketCore.scala 283:16]
  wire  _T_872; // @[RocketCore.scala 282:48]
  wire  _T_875; // @[RocketCore.scala 284:16]
  wire  _T_876; // @[RocketCore.scala 283:70]
  wire  _T_879; // @[RocketCore.scala 285:30]
  wire  _T_880; // @[RocketCore.scala 284:47]
  wire  _T_886; // @[RocketCore.scala 288:64]
  wire  _T_887; // @[RocketCore.scala 288:49]
  wire  _T_888; // @[RocketCore.scala 288:15]
  wire  _T_889; // @[RocketCore.scala 287:73]
  wire  _T_892; // @[RocketCore.scala 289:65]
  wire  _T_893; // @[RocketCore.scala 289:31]
  wire  id_illegal_insn; // @[RocketCore.scala 288:99]
  wire  id_amo_aq; // @[RocketCore.scala 291:29]
  wire  id_amo_rl; // @[RocketCore.scala 292:29]
  wire  _T_894; // @[RocketCore.scala 293:52]
  wire  id_fence_next; // @[RocketCore.scala 293:37]
  wire  id_mem_busy; // @[RocketCore.scala 294:38]
  wire  _GEN_0; // @[RocketCore.scala 295:23]
  wire  _T_904; // @[RocketCore.scala 300:33]
  wire  _T_905; // @[RocketCore.scala 300:46]
  wire  _T_907; // @[RocketCore.scala 300:81]
  wire  _T_908; // @[RocketCore.scala 300:65]
  wire  id_do_fence; // @[RocketCore.scala 300:17]
  wire  _T_912; // @[RocketCore.scala 892:26]
  wire  _T_913; // @[RocketCore.scala 892:26]
  wire  _T_914; // @[RocketCore.scala 892:26]
  wire  _T_915; // @[RocketCore.scala 892:26]
  wire  _T_916; // @[RocketCore.scala 892:26]
  wire  _T_917; // @[RocketCore.scala 892:26]
  wire  id_xcpt; // @[RocketCore.scala 892:26]
  wire [1:0] _T_918; // @[Mux.scala 31:69]
  wire [3:0] _T_919; // @[Mux.scala 31:69]
  wire [3:0] _T_920; // @[Mux.scala 31:69]
  wire [3:0] _T_921; // @[Mux.scala 31:69]
  wire [3:0] _T_922; // @[Mux.scala 31:69]
  wire [3:0] _T_923; // @[Mux.scala 31:69]
  wire [4:0] ex_waddr; // @[RocketCore.scala 335:29]
  wire [4:0] mem_waddr; // @[RocketCore.scala 336:31]
  wire [4:0] wb_waddr; // @[RocketCore.scala 337:29]
  wire  _T_934; // @[RocketCore.scala 340:19]
  wire  _T_935; // @[RocketCore.scala 341:20]
  wire  _T_937; // @[RocketCore.scala 341:36]
  wire  _T_939; // @[RocketCore.scala 343:82]
  wire  _T_941; // @[RocketCore.scala 343:82]
  wire  _T_942; // @[RocketCore.scala 343:74]
  wire  _T_943; // @[RocketCore.scala 343:82]
  wire  _T_944; // @[RocketCore.scala 343:74]
  wire  _T_946; // @[RocketCore.scala 343:74]
  wire  _T_947; // @[RocketCore.scala 343:82]
  wire  _T_949; // @[RocketCore.scala 343:82]
  wire  _T_950; // @[RocketCore.scala 343:74]
  wire  _T_951; // @[RocketCore.scala 343:82]
  wire  _T_952; // @[RocketCore.scala 343:74]
  wire  _T_954; // @[RocketCore.scala 343:74]
  reg  ex_reg_rs_bypass_0; // @[RocketCore.scala 347:29]
  reg [31:0] _RAND_80;
  reg  ex_reg_rs_bypass_1; // @[RocketCore.scala 347:29]
  reg [31:0] _RAND_81;
  reg [1:0] ex_reg_rs_lsb_0; // @[RocketCore.scala 348:26]
  reg [31:0] _RAND_82;
  reg [1:0] ex_reg_rs_lsb_1; // @[RocketCore.scala 348:26]
  reg [31:0] _RAND_83;
  reg [61:0] ex_reg_rs_msb_0; // @[RocketCore.scala 349:26]
  reg [63:0] _RAND_84;
  reg [61:0] ex_reg_rs_msb_1; // @[RocketCore.scala 349:26]
  reg [63:0] _RAND_85;
  wire  _T_976; // @[package.scala 31:81]
  wire [63:0] _T_977; // @[package.scala 31:71]
  wire  _T_978; // @[package.scala 31:81]
  wire [63:0] _T_979; // @[package.scala 31:71]
  wire  _T_980; // @[package.scala 31:81]
  wire [63:0] _T_981; // @[package.scala 31:71]
  wire [63:0] _T_982; // @[Cat.scala 30:58]
  wire  _T_984; // @[package.scala 31:81]
  wire [63:0] _T_985; // @[package.scala 31:71]
  wire  _T_986; // @[package.scala 31:81]
  wire [63:0] _T_987; // @[package.scala 31:71]
  wire  _T_988; // @[package.scala 31:81]
  wire [63:0] _T_989; // @[package.scala 31:71]
  wire [63:0] _T_990; // @[Cat.scala 30:58]
  wire [63:0] _T_991; // @[RocketCore.scala 351:14]
  wire  _T_992; // @[RocketCore.scala 954:24]
  wire  _T_994; // @[RocketCore.scala 954:53]
  wire  _T_995; // @[RocketCore.scala 954:19]
  wire  _T_996; // @[RocketCore.scala 955:26]
  wire [10:0] _T_998; // @[RocketCore.scala 955:49]
  wire  _T_1000; // @[RocketCore.scala 956:26]
  wire  _T_1001; // @[RocketCore.scala 956:43]
  wire  _T_1002; // @[RocketCore.scala 956:36]
  wire [7:0] _T_1004; // @[RocketCore.scala 956:73]
  wire  _T_1008; // @[RocketCore.scala 957:33]
  wire  _T_1009; // @[RocketCore.scala 958:23]
  wire  _T_1011; // @[RocketCore.scala 958:44]
  wire  _T_1012; // @[RocketCore.scala 959:23]
  wire  _T_1014; // @[RocketCore.scala 959:43]
  wire  _T_1015; // @[RocketCore.scala 959:18]
  wire  _T_1016; // @[RocketCore.scala 958:18]
  wire [5:0] _T_1022; // @[RocketCore.scala 960:20]
  wire  _T_1024; // @[RocketCore.scala 962:24]
  wire  _T_1026; // @[RocketCore.scala 962:34]
  wire [3:0] _T_1031; // @[RocketCore.scala 963:19]
  wire [3:0] _T_1032; // @[RocketCore.scala 962:19]
  wire [3:0] _T_1033; // @[RocketCore.scala 961:19]
  wire  _T_1036; // @[RocketCore.scala 965:22]
  wire  _T_1040; // @[RocketCore.scala 966:17]
  wire  _T_1041; // @[RocketCore.scala 965:17]
  wire  _T_1042; // @[RocketCore.scala 964:17]
  wire  _T_1045; // @[Cat.scala 30:58]
  wire [7:0] _T_1046; // @[Cat.scala 30:58]
  wire [10:0] _T_1048; // @[Cat.scala 30:58]
  wire  _T_1049; // @[Cat.scala 30:58]
  wire [31:0] ex_imm; // @[RocketCore.scala 968:53]
  wire [63:0] _T_1053; // @[RocketCore.scala 354:24]
  wire  _T_1055; // @[Mux.scala 46:19]
  wire [39:0] _T_1056; // @[Mux.scala 46:16]
  wire  _T_1057; // @[Mux.scala 46:19]
  wire [63:0] _T_1058; // @[RocketCore.scala 357:24]
  wire [3:0] _T_1059; // @[RocketCore.scala 359:19]
  wire  _T_1060; // @[Mux.scala 46:19]
  wire [3:0] _T_1061; // @[Mux.scala 46:16]
  wire  _T_1062; // @[Mux.scala 46:19]
  wire [31:0] _T_1063; // @[Mux.scala 46:16]
  wire  _T_1064; // @[Mux.scala 46:19]
  wire  _T_1739; // @[RocketCore.scala 724:40]
  wire  _T_1740; // @[RocketCore.scala 724:71]
  wire  _T_1543; // @[RocketCore.scala 656:55]
  wire  _T_1544; // @[RocketCore.scala 656:42]
  wire  _T_1591; // @[RocketCore.scala 676:70]
  wire  _T_1592; // @[RocketCore.scala 901:27]
  wire  _T_1545; // @[RocketCore.scala 657:55]
  wire  _T_1546; // @[RocketCore.scala 657:42]
  wire  _T_1593; // @[RocketCore.scala 676:70]
  wire  _T_1594; // @[RocketCore.scala 901:27]
  wire  _T_1597; // @[RocketCore.scala 901:50]
  wire  _T_1547; // @[RocketCore.scala 658:55]
  wire  _T_1548; // @[RocketCore.scala 658:42]
  wire  _T_1595; // @[RocketCore.scala 676:70]
  wire  _T_1596; // @[RocketCore.scala 901:27]
  wire  _T_1598; // @[RocketCore.scala 901:50]
  wire  data_hazard_ex; // @[RocketCore.scala 676:36]
  wire  _T_1585; // @[RocketCore.scala 675:38]
  wire  _T_1586; // @[RocketCore.scala 675:48]
  wire  _T_1587; // @[RocketCore.scala 675:64]
  wire  _T_1589; // @[RocketCore.scala 675:94]
  wire  ex_cannot_bypass; // @[RocketCore.scala 675:109]
  wire  _T_1610; // @[RocketCore.scala 678:54]
  wire  _T_1600; // @[RocketCore.scala 901:27]
  wire  _T_1602; // @[RocketCore.scala 901:27]
  wire  _T_1607; // @[RocketCore.scala 901:50]
  wire  _T_1603; // @[RocketCore.scala 677:76]
  wire  _T_1604; // @[RocketCore.scala 901:27]
  wire  _T_1608; // @[RocketCore.scala 901:50]
  wire  _T_1606; // @[RocketCore.scala 901:27]
  wire  _T_1609; // @[RocketCore.scala 901:50]
  wire  fp_data_hazard_ex; // @[RocketCore.scala 677:39]
  wire  _T_1611; // @[RocketCore.scala 678:74]
  wire  id_ex_hazard; // @[RocketCore.scala 678:35]
  wire  _T_1618; // @[RocketCore.scala 685:72]
  wire  _T_1619; // @[RocketCore.scala 901:27]
  wire  _T_1620; // @[RocketCore.scala 685:72]
  wire  _T_1621; // @[RocketCore.scala 901:27]
  wire  _T_1624; // @[RocketCore.scala 901:50]
  wire  _T_1622; // @[RocketCore.scala 685:72]
  wire  _T_1623; // @[RocketCore.scala 901:27]
  wire  _T_1625; // @[RocketCore.scala 901:50]
  wire  data_hazard_mem; // @[RocketCore.scala 685:38]
  wire  _T_1612; // @[RocketCore.scala 684:40]
  wire  _T_1613; // @[RocketCore.scala 684:66]
  wire  _T_1614; // @[RocketCore.scala 684:50]
  wire  _T_1616; // @[RocketCore.scala 684:100]
  wire  mem_cannot_bypass; // @[RocketCore.scala 684:116]
  wire  _T_1637; // @[RocketCore.scala 687:57]
  wire  _T_1627; // @[RocketCore.scala 901:27]
  wire  _T_1629; // @[RocketCore.scala 901:27]
  wire  _T_1634; // @[RocketCore.scala 901:50]
  wire  _T_1630; // @[RocketCore.scala 686:78]
  wire  _T_1631; // @[RocketCore.scala 901:27]
  wire  _T_1635; // @[RocketCore.scala 901:50]
  wire  _T_1633; // @[RocketCore.scala 901:27]
  wire  _T_1636; // @[RocketCore.scala 901:50]
  wire  fp_data_hazard_mem; // @[RocketCore.scala 686:41]
  wire  _T_1638; // @[RocketCore.scala 687:78]
  wire  id_mem_hazard; // @[RocketCore.scala 687:37]
  wire  _T_1711; // @[RocketCore.scala 714:18]
  wire  _T_1641; // @[RocketCore.scala 691:70]
  wire  _T_1642; // @[RocketCore.scala 901:27]
  wire  _T_1643; // @[RocketCore.scala 691:70]
  wire  _T_1644; // @[RocketCore.scala 901:27]
  wire  _T_1647; // @[RocketCore.scala 901:50]
  wire  _T_1645; // @[RocketCore.scala 691:70]
  wire  _T_1646; // @[RocketCore.scala 901:27]
  wire  _T_1648; // @[RocketCore.scala 901:50]
  wire  data_hazard_wb; // @[RocketCore.scala 691:36]
  wire  wb_dcache_miss; // @[RocketCore.scala 448:36]
  wire  wb_set_sboard; // @[RocketCore.scala 584:35]
  wire  _T_1660; // @[RocketCore.scala 693:54]
  wire  _T_1650; // @[RocketCore.scala 901:27]
  wire  _T_1652; // @[RocketCore.scala 901:27]
  wire  _T_1657; // @[RocketCore.scala 901:50]
  wire  _T_1653; // @[RocketCore.scala 692:76]
  wire  _T_1654; // @[RocketCore.scala 901:27]
  wire  _T_1658; // @[RocketCore.scala 901:50]
  wire  _T_1656; // @[RocketCore.scala 901:27]
  wire  _T_1659; // @[RocketCore.scala 901:50]
  wire  fp_data_hazard_wb; // @[RocketCore.scala 692:39]
  wire  _T_1661; // @[RocketCore.scala 693:71]
  wire  id_wb_hazard; // @[RocketCore.scala 693:35]
  wire  _T_1712; // @[RocketCore.scala 714:35]
  reg [31:0] _T_1550; // @[RocketCore.scala 918:25]
  reg [31:0] _RAND_86;
  wire [31:0] _T_1552; // @[RocketCore.scala 919:40]
  wire [31:0] _T_1558; // @[RocketCore.scala 915:35]
  wire  dmem_resp_valid; // @[RocketCore.scala 594:44]
  wire  dmem_resp_replay; // @[RocketCore.scala 595:42]
  wire  dmem_resp_xpu; // @[RocketCore.scala 591:23]
  wire  _T_1486; // @[RocketCore.scala 610:26]
  wire  _T_1484; // @[Decoupled.scala 37:37]
  wire  ll_wen; // @[RocketCore.scala 610:44]
  wire [4:0] dmem_resp_waddr; // @[RocketCore.scala 593:46]
  wire [4:0] ll_waddr; // @[RocketCore.scala 610:44]
  wire  _T_1560; // @[RocketCore.scala 668:70]
  wire  _T_1561; // @[RocketCore.scala 668:58]
  wire  _T_1563; // @[RocketCore.scala 671:77]
  wire  _T_1564; // @[RocketCore.scala 901:27]
  wire [31:0] _T_1565; // @[RocketCore.scala 915:35]
  wire  _T_1567; // @[RocketCore.scala 668:70]
  wire  _T_1568; // @[RocketCore.scala 668:58]
  wire  _T_1570; // @[RocketCore.scala 671:77]
  wire  _T_1571; // @[RocketCore.scala 901:27]
  wire  _T_1579; // @[RocketCore.scala 901:50]
  wire [31:0] _T_1572; // @[RocketCore.scala 915:35]
  wire  _T_1574; // @[RocketCore.scala 668:70]
  wire  _T_1575; // @[RocketCore.scala 668:58]
  wire  _T_1577; // @[RocketCore.scala 671:77]
  wire  _T_1578; // @[RocketCore.scala 901:27]
  wire  id_sboard_hazard; // @[RocketCore.scala 901:50]
  wire  _T_1713; // @[RocketCore.scala 714:51]
  wire  _T_1714; // @[RocketCore.scala 715:40]
  wire  _T_1715; // @[RocketCore.scala 715:57]
  wire  _T_1716; // @[RocketCore.scala 715:23]
  wire  _T_1717; // @[RocketCore.scala 714:71]
  wire  _T_1718; // @[RocketCore.scala 716:15]
  wire  _T_1720; // @[RocketCore.scala 716:42]
  wire  _T_1721; // @[RocketCore.scala 715:74]
  reg [31:0] _T_1663; // @[RocketCore.scala 918:25]
  reg [31:0] _RAND_87;
  wire [31:0] _T_1682; // @[RocketCore.scala 915:35]
  wire  _T_1684; // @[RocketCore.scala 901:27]
  wire [31:0] _T_1685; // @[RocketCore.scala 915:35]
  wire  _T_1687; // @[RocketCore.scala 901:27]
  wire  _T_1694; // @[RocketCore.scala 901:50]
  wire [31:0] _T_1688; // @[RocketCore.scala 915:35]
  wire  _T_1690; // @[RocketCore.scala 901:27]
  wire  _T_1695; // @[RocketCore.scala 901:50]
  wire [31:0] _T_1691; // @[RocketCore.scala 915:35]
  wire  _T_1693; // @[RocketCore.scala 901:27]
  wire  id_stall_fpu; // @[RocketCore.scala 901:50]
  wire  _T_1722; // @[RocketCore.scala 717:16]
  wire  _T_1723; // @[RocketCore.scala 716:62]
  reg  blocked; // @[RocketCore.scala 706:22]
  reg [31:0] _RAND_88;
  wire  dcache_blocked; // @[RocketCore.scala 708:13]
  wire  _T_1724; // @[RocketCore.scala 718:17]
  wire  _T_1725; // @[RocketCore.scala 717:32]
  wire  wb_wxd; // @[RocketCore.scala 583:29]
  wire  _T_1729; // @[RocketCore.scala 720:62]
  wire  _T_1730; // @[RocketCore.scala 720:40]
  wire  _T_1732; // @[RocketCore.scala 720:75]
  wire  _T_1733; // @[RocketCore.scala 720:17]
  wire  _T_1734; // @[RocketCore.scala 719:34]
  wire  _T_1737; // @[RocketCore.scala 721:15]
  wire  ctrl_stalld; // @[RocketCore.scala 722:17]
  wire  _T_1741; // @[RocketCore.scala 724:89]
  wire  ctrl_killd; // @[RocketCore.scala 724:104]
  wire  _T_1070; // @[RocketCore.scala 391:29]
  wire  _GEN_1; // @[RocketCore.scala 399:26]
  wire [1:0] _T_1078; // @[RocketCore.scala 405:22]
  wire  _T_1079; // @[RocketCore.scala 405:29]
  wire  _GEN_4; // @[RocketCore.scala 405:34]
  wire [1:0] _T_1080; // @[RocketCore.scala 410:40]
  wire  _T_1081; // @[RocketCore.scala 410:47]
  wire  _T_1082; // @[RocketCore.scala 410:28]
  wire  _GEN_8; // @[RocketCore.scala 400:20]
  wire  _T_1083; // @[RocketCore.scala 415:42]
  wire [1:0] _T_1086; // @[Cat.scala 30:58]
  wire  _T_1087; // @[RocketCore.scala 422:48]
  wire  _T_1088; // @[RocketCore.scala 422:48]
  wire  do_bypass; // @[RocketCore.scala 422:48]
  wire  _T_1092; // @[RocketCore.scala 426:23]
  wire  _T_1488; // @[RocketCore.scala 618:31]
  wire  wb_valid; // @[RocketCore.scala 618:45]
  wire  wb_wen; // @[RocketCore.scala 619:25]
  wire  rf_wen; // @[RocketCore.scala 620:23]
  wire [4:0] rf_waddr; // @[RocketCore.scala 621:21]
  wire  _T_1496; // @[RocketCore.scala 944:16]
  wire  _T_1500; // @[RocketCore.scala 947:20]
  wire  _T_1490; // @[RocketCore.scala 622:38]
  wire [63:0] ll_wdata;
  wire  _T_1492; // @[RocketCore.scala 624:34]
  wire [63:0] _T_1494; // @[RocketCore.scala 624:21]
  wire [63:0] _T_1495; // @[RocketCore.scala 623:21]
  wire [63:0] rf_wdata; // @[RocketCore.scala 622:21]
  wire [63:0] _GEN_214; // @[RocketCore.scala 947:31]
  wire [63:0] _GEN_221; // @[RocketCore.scala 944:29]
  wire [63:0] _GEN_228; // @[RocketCore.scala 627:17]
  wire  _T_1095; // @[RocketCore.scala 422:48]
  wire  _T_1096; // @[RocketCore.scala 422:48]
  wire  do_bypass_1; // @[RocketCore.scala 422:48]
  wire  _T_1100; // @[RocketCore.scala 426:23]
  wire  _T_1501; // @[RocketCore.scala 947:20]
  wire [63:0] _GEN_215; // @[RocketCore.scala 947:31]
  wire [63:0] _GEN_222; // @[RocketCore.scala 944:29]
  wire [63:0] _GEN_229; // @[RocketCore.scala 627:17]
  wire [31:0] inst; // @[RocketCore.scala 432:21]
  wire  _T_1639; // @[RocketCore.scala 688:32]
  wire  id_load_use; // @[RocketCore.scala 688:51]
  wire  _T_1107; // @[RocketCore.scala 438:21]
  wire  _T_1108; // @[RocketCore.scala 438:41]
  wire  _T_1112; // @[RocketCore.scala 449:42]
  wire  _T_1114; // @[RocketCore.scala 450:42]
  wire  replay_ex_structural; // @[RocketCore.scala 449:64]
  wire  replay_ex_load_use; // @[RocketCore.scala 451:43]
  wire  _T_1115; // @[RocketCore.scala 452:75]
  wire  _T_1116; // @[RocketCore.scala 452:50]
  wire  replay_ex; // @[RocketCore.scala 452:33]
  wire  _T_1117; // @[RocketCore.scala 453:35]
  wire  ctrl_killx; // @[RocketCore.scala 453:48]
  wire  _T_1119; // @[RocketCore.scala 455:40]
  wire  _T_1130; // @[RocketCore.scala 455:91]
  wire  _T_1131; // @[RocketCore.scala 455:91]
  wire  _T_1132; // @[RocketCore.scala 455:91]
  wire  _T_1133; // @[RocketCore.scala 455:91]
  wire  _T_1135; // @[RocketCore.scala 455:91]
  wire  _T_1136; // @[RocketCore.scala 455:91]
  wire  _T_1137; // @[RocketCore.scala 455:91]
  wire  ex_slow_bypass; // @[RocketCore.scala 455:50]
  wire  _T_1139; // @[RocketCore.scala 456:67]
  wire  ex_sfence; // @[RocketCore.scala 456:48]
  wire  ex_xcpt; // @[RocketCore.scala 459:28]
  wire  _T_1150; // @[RocketCore.scala 465:36]
  wire  mem_pc_valid; // @[RocketCore.scala 465:54]
  wire  _T_1303; // @[RocketCore.scala 474:56]
  wire  mem_npc_misaligned; // @[RocketCore.scala 474:70]
  wire  _T_1306; // @[RocketCore.scala 475:59]
  wire  _T_1307; // @[RocketCore.scala 475:41]
  wire [63:0] mem_int_wdata; // @[RocketCore.scala 475:119]
  wire  _T_1310; // @[RocketCore.scala 476:33]
  wire  mem_cfi; // @[RocketCore.scala 476:50]
  wire  _T_1312; // @[RocketCore.scala 477:57]
  wire  mem_cfi_taken; // @[RocketCore.scala 477:74]
  wire  _T_1324; // @[RocketCore.scala 489:23]
  wire  _T_1325; // @[Consts.scala 93:31]
  wire  _T_1326; // @[Consts.scala 93:48]
  wire  _T_1327; // @[Consts.scala 93:41]
  wire  _T_1329; // @[Consts.scala 93:58]
  wire  _T_1330; // @[package.scala 14:47]
  wire  _T_1331; // @[package.scala 14:47]
  wire  _T_1332; // @[package.scala 14:47]
  wire  _T_1333; // @[package.scala 14:47]
  wire  _T_1334; // @[package.scala 14:62]
  wire  _T_1335; // @[package.scala 14:62]
  wire  _T_1336; // @[package.scala 14:62]
  wire  _T_1337; // @[package.scala 14:47]
  wire  _T_1338; // @[package.scala 14:47]
  wire  _T_1339; // @[package.scala 14:47]
  wire  _T_1340; // @[package.scala 14:47]
  wire  _T_1341; // @[package.scala 14:47]
  wire  _T_1342; // @[package.scala 14:62]
  wire  _T_1343; // @[package.scala 14:62]
  wire  _T_1344; // @[package.scala 14:62]
  wire  _T_1345; // @[package.scala 14:62]
  wire  _T_1346; // @[Consts.scala 91:44]
  wire  _T_1347; // @[Consts.scala 93:75]
  wire  _T_1348; // @[RocketCore.scala 494:33]
  wire  _T_1349; // @[Consts.scala 94:32]
  wire  _T_1350; // @[Consts.scala 94:49]
  wire  _T_1351; // @[Consts.scala 94:42]
  wire  _T_1353; // @[Consts.scala 94:59]
  wire  _T_1371; // @[Consts.scala 94:76]
  wire  _T_1372; // @[RocketCore.scala 495:34]
  wire  _T_1374; // @[RocketCore.scala 508:56]
  wire  _T_1375; // @[RocketCore.scala 508:24]
  wire  _T_1377; // @[AMOALU.scala 26:19]
  wire [63:0] _T_1381; // @[Cat.scala 30:58]
  wire  _T_1382; // @[AMOALU.scala 26:19]
  wire [63:0] _T_1385; // @[Cat.scala 30:58]
  wire  _T_1386; // @[AMOALU.scala 26:19]
  wire [63:0] _T_1388; // @[Cat.scala 30:58]
  wire  _T_1392; // @[RocketCore.scala 512:24]
  wire  _GEN_72; // @[RocketCore.scala 512:48]
  wire  _GEN_73; // @[RocketCore.scala 512:48]
  wire  _T_1393; // @[RocketCore.scala 519:38]
  wire  _T_1394; // @[RocketCore.scala 519:75]
  wire  mem_breakpoint; // @[RocketCore.scala 519:57]
  wire  _T_1395; // @[RocketCore.scala 520:44]
  wire  _T_1396; // @[RocketCore.scala 520:82]
  wire  mem_debug_breakpoint; // @[RocketCore.scala 520:64]
  wire  mem_ldst_xcpt; // @[RocketCore.scala 892:26]
  wire [3:0] mem_ldst_cause; // @[Mux.scala 31:69]
  wire  _T_1397; // @[RocketCore.scala 526:29]
  wire  _T_1398; // @[RocketCore.scala 527:20]
  wire  _T_1399; // @[RocketCore.scala 528:20]
  wire  _T_1400; // @[RocketCore.scala 892:26]
  wire  mem_xcpt; // @[RocketCore.scala 892:26]
  wire [3:0] _T_1401; // @[Mux.scala 31:69]
  wire  dcache_kill_mem; // @[RocketCore.scala 537:55]
  wire  _T_1415; // @[RocketCore.scala 538:36]
  wire  fpu_kill_mem; // @[RocketCore.scala 538:51]
  wire  _T_1416; // @[RocketCore.scala 539:37]
  wire  replay_mem; // @[RocketCore.scala 539:55]
  wire  _T_1417; // @[RocketCore.scala 540:38]
  wire  _T_1418; // @[RocketCore.scala 540:52]
  wire  killm_common; // @[RocketCore.scala 540:68]
  reg  _T_1422; // @[RocketCore.scala 541:37]
  reg [31:0] _RAND_89;
  wire  _T_1424; // @[RocketCore.scala 542:33]
  wire  ctrl_killm; // @[RocketCore.scala 542:45]
  wire  _T_1433; // @[RocketCore.scala 552:39]
  wire  _T_1434; // @[RocketCore.scala 552:54]
  wire [2:0] _T_1454; // @[Mux.scala 31:69]
  wire [3:0] _T_1455; // @[Mux.scala 31:69]
  wire [3:0] _T_1456; // @[Mux.scala 31:69]
  wire [3:0] _T_1457; // @[Mux.scala 31:69]
  wire [3:0] _T_1458; // @[Mux.scala 31:69]
  wire [63:0] wb_cause; // @[Mux.scala 31:69]
  wire  _T_1459; // @[RocketCore.scala 896:38]
  wire  _T_1461; // @[RocketCore.scala 896:38]
  wire  _T_1463; // @[RocketCore.scala 896:38]
  wire  _T_1465; // @[RocketCore.scala 896:38]
  wire  _T_1467; // @[RocketCore.scala 896:38]
  wire  _T_1469; // @[RocketCore.scala 896:38]
  wire  _T_1510; // @[package.scala 14:47]
  wire  _T_1511; // @[package.scala 14:47]
  wire  _T_1516; // @[package.scala 14:47]
  wire  _T_1519; // @[package.scala 14:47]
  wire  _T_1520; // @[package.scala 14:62]
  wire  _T_1521; // @[package.scala 14:62]
  wire  _T_1522; // @[package.scala 14:62]
  wire  _T_1523; // @[package.scala 14:62]
  wire  _T_1524; // @[package.scala 14:62]
  wire  _T_1525; // @[package.scala 14:62]
  wire  _T_1526; // @[package.scala 14:62]
  wire  _T_1527; // @[package.scala 14:62]
  wire  _T_1528; // @[package.scala 14:62]
  wire  tval_valid; // @[RocketCore.scala 642:28]
  wire [24:0] a_1; // @[RocketCore.scala 906:23]
  wire  _T_1530; // @[RocketCore.scala 907:21]
  wire  _T_1531; // @[RocketCore.scala 907:34]
  wire  _T_1532; // @[RocketCore.scala 907:29]
  wire  msb_1; // @[RocketCore.scala 907:18]
  wire [39:0] _T_1537; // @[Cat.scala 30:58]
  wire [2:0] _T_1540; // @[CSR.scala 128:15]
  wire [31:0] _T_1553; // @[RocketCore.scala 922:62]
  wire [31:0] _T_1554; // @[RocketCore.scala 922:49]
  wire [31:0] _T_1556; // @[RocketCore.scala 914:62]
  wire  _T_1580; // @[RocketCore.scala 672:28]
  wire [31:0] _T_1581; // @[RocketCore.scala 922:62]
  wire [31:0] _T_1582; // @[RocketCore.scala 922:49]
  wire [31:0] _T_1583; // @[RocketCore.scala 913:60]
  wire  _T_1584; // @[RocketCore.scala 925:17]
  wire  _T_1664; // @[RocketCore.scala 697:35]
  wire  _T_1665; // @[RocketCore.scala 697:50]
  wire  _T_1666; // @[RocketCore.scala 697:72]
  wire [31:0] _T_1668; // @[RocketCore.scala 922:49]
  wire [31:0] _T_1669; // @[RocketCore.scala 913:60]
  wire  _T_1671; // @[RocketCore.scala 698:38]
  wire [31:0] _T_1672; // @[RocketCore.scala 922:62]
  wire [31:0] _T_1673; // @[RocketCore.scala 922:49]
  wire [31:0] _T_1675; // @[RocketCore.scala 914:62]
  wire  _T_1676; // @[RocketCore.scala 925:17]
  wire [31:0] _T_1677; // @[RocketCore.scala 922:62]
  wire [31:0] _T_1678; // @[RocketCore.scala 922:49]
  wire [31:0] _T_1680; // @[RocketCore.scala 914:62]
  wire  _T_1681; // @[RocketCore.scala 925:17]
  wire  _T_1698; // @[RocketCore.scala 707:35]
  wire  _T_1700; // @[RocketCore.scala 707:60]
  wire  _T_1701; // @[RocketCore.scala 707:95]
  wire  _T_1702; // @[RocketCore.scala 707:116]
  wire  _T_1744; // @[RocketCore.scala 729:17]
  wire [39:0] _T_1745; // @[RocketCore.scala 730:8]
  wire  _T_1747; // @[RocketCore.scala 732:40]
  wire  _T_1750; // @[RocketCore.scala 734:43]
  wire  _T_1758; // @[RocketCore.scala 746:45]
  wire  _T_1759; // @[RocketCore.scala 746:60]
  wire  _T_1761; // @[RocketCore.scala 746:90]
  wire  _T_1763; // @[RocketCore.scala 749:23]
  wire  _T_1765; // @[RocketCore.scala 749:41]
  wire [4:0] _T_1767; // @[RocketCore.scala 750:46]
  wire  _T_1768; // @[RocketCore.scala 750:46]
  wire  _T_1769; // @[RocketCore.scala 750:23]
  wire [1:0] _T_1772; // @[RocketCore.scala 750:8]
  wire [1:0] _T_1774; // @[RocketCore.scala 754:74]
  wire [39:0] _GEN_237; // @[RocketCore.scala 754:69]
  wire [39:0] _T_1776; // @[RocketCore.scala 754:69]
  wire [38:0] _T_1778; // @[RocketCore.scala 755:66]
  wire [5:0] ex_dcache_tag; // @[Cat.scala 30:58]
  wire [24:0] a_2; // @[RocketCore.scala 906:23]
  wire  _T_1788; // @[RocketCore.scala 907:21]
  wire  _T_1789; // @[RocketCore.scala 907:34]
  wire  _T_1790; // @[RocketCore.scala 907:29]
  wire  msb_2; // @[RocketCore.scala 907:18]
  wire  _T_1797; // @[RocketCore.scala 785:35]
  reg [19:0] Rocket_state; // @[Register tracking Rocket state]
  reg [31:0] _RAND_90;
  reg  Rocket_cov [0:1048575]; // @[Coverage map for Rocket]
  reg [31:0] _RAND_91;
  wire  Rocket_cov_read_data; // @[Coverage map for Rocket]
  wire [19:0] Rocket_cov_read_addr; // @[Coverage map for Rocket]
  wire  Rocket_cov_write_data; // @[Coverage map for Rocket]
  wire [19:0] Rocket_cov_write_addr; // @[Coverage map for Rocket]
  wire  Rocket_cov_write_mask; // @[Coverage map for Rocket]
  wire  Rocket_cov_write_en; // @[Coverage map for Rocket]
  reg [29:0] Rocket_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_92;
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  mux_cond_4;
  wire [1:0] wb_ctrl_wfd_shl;
  wire [19:0] wb_ctrl_wfd_pad;
  wire [6:0] ex_ctrl_mem_type_shl;
  wire [19:0] ex_ctrl_mem_type_pad;
  wire [8:0] wb_reg_replay_shl;
  wire [19:0] wb_reg_replay_pad;
  wire [19:0] wb_ctrl_mem_shl;
  wire [19:0] wb_ctrl_mem_pad;
  wire [11:0] mem_ctrl_jalr_shl;
  wire [19:0] mem_ctrl_jalr_pad;
  wire [3:0] ex_ctrl_wfd_shl;
  wire [19:0] ex_ctrl_wfd_pad;
  wire [1:0] mem_ctrl_wfd_shl;
  wire [19:0] mem_ctrl_wfd_pad;
  wire [15:0] ex_ctrl_sel_alu1_shl;
  wire [19:0] ex_ctrl_sel_alu1_pad;
  wire [19:0] ex_ctrl_fp_shl;
  wire [19:0] ex_ctrl_fp_pad;
  wire [2:0] mem_reg_rvc_shl;
  wire [19:0] mem_reg_rvc_pad;
  wire [5:0] ex_ctrl_rxs2_shl;
  wire [19:0] ex_ctrl_rxs2_pad;
  wire [3:0] ex_reg_xcpt_interrupt_shl;
  wire [19:0] ex_reg_xcpt_interrupt_pad;
  wire [4:0] mem_reg_valid_shl;
  wire [19:0] mem_reg_valid_pad;
  wire [6:0] mem_ctrl_mem_shl;
  wire [19:0] mem_ctrl_mem_pad;
  wire  mem_reg_store_shl;
  wire [19:0] mem_reg_store_pad;
  wire [6:0] mem_reg_xcpt_shl;
  wire [19:0] mem_reg_xcpt_pad;
  wire [1:0] mem_ctrl_branch_shl;
  wire [19:0] mem_ctrl_branch_pad;
  wire [11:0] ex_ctrl_wxd_shl;
  wire [19:0] ex_ctrl_wxd_pad;
  wire [2:0] mem_ctrl_wxd_shl;
  wire [19:0] mem_ctrl_wxd_pad;
  wire [7:0] ex_ctrl_mem_shl;
  wire [19:0] ex_ctrl_mem_pad;
  wire [3:0] mem_reg_replay_shl;
  wire [19:0] mem_reg_replay_pad;
  wire [8:0] wb_reg_xcpt_shl;
  wire [19:0] wb_reg_xcpt_pad;
  wire [9:0] mem_ctrl_jal_shl;
  wire [19:0] mem_ctrl_jal_pad;
  wire [1:0] ex_ctrl_jalr_shl;
  wire [19:0] ex_ctrl_jalr_pad;
  wire [17:0] mem_reg_flush_pipe_shl;
  wire [19:0] mem_reg_flush_pipe_pad;
  wire [10:0] mem_reg_xcpt_interrupt_shl;
  wire [19:0] mem_reg_xcpt_interrupt_pad;
  wire [7:0] ex_reg_replay_shl;
  wire [19:0] ex_reg_replay_pad;
  wire [13:0] ex_ctrl_sel_alu2_shl;
  wire [19:0] ex_ctrl_sel_alu2_pad;
  wire [5:0] ex_reg_valid_shl;
  wire [19:0] ex_reg_valid_pad;
  wire [9:0] mem_ctrl_fp_shl;
  wire [19:0] mem_ctrl_fp_pad;
  wire [12:0] id_reg_fence_shl;
  wire [19:0] id_reg_fence_pad;
  wire [1:0] wb_ctrl_div_shl;
  wire [19:0] wb_ctrl_div_pad;
  wire [4:0] ex_ctrl_sel_imm_shl;
  wire [19:0] ex_ctrl_sel_imm_pad;
  wire [9:0] wb_ctrl_wxd_shl;
  wire [19:0] wb_ctrl_wxd_pad;
  wire [12:0] ex_ctrl_div_shl;
  wire [19:0] ex_ctrl_div_pad;
  wire [14:0] wb_reg_valid_shl;
  wire [19:0] wb_reg_valid_pad;
  wire [9:0] mem_reg_sfence_shl;
  wire [19:0] mem_reg_sfence_pad;
  wire [9:0] ex_reg_rvc_shl;
  wire [19:0] ex_reg_rvc_pad;
  wire [19:0] mem_reg_load_shl;
  wire [19:0] mem_reg_load_pad;
  wire [13:0] wb_reg_flush_pipe_shl;
  wire [19:0] wb_reg_flush_pipe_pad;
  wire [10:0] mem_reg_slow_bypass_shl;
  wire [19:0] mem_reg_slow_bypass_pad;
  wire [8:0] blocked_shl;
  wire [19:0] blocked_pad;
  wire [9:0] mem_br_taken_shl;
  wire [19:0] mem_br_taken_pad;
  wire [6:0] mem_ctrl_div_shl;
  wire [19:0] mem_ctrl_div_pad;
  wire [13:0] mux_cond_0_shl;
  wire [19:0] mux_cond_0_pad;
  wire [15:0] mux_cond_1_shl;
  wire [19:0] mux_cond_1_pad;
  wire [7:0] mux_cond_2_shl;
  wire [19:0] mux_cond_2_pad;
  wire [8:0] mux_cond_3_shl;
  wire [19:0] mux_cond_3_pad;
  wire [1:0] mux_cond_4_shl;
  wire [19:0] mux_cond_4_pad;
  wire [8:0] ex_reg_rs_bypass_0_shl;
  wire [19:0] ex_reg_rs_bypass_0_pad;
  wire [8:0] ex_reg_rs_bypass_1_shl;
  wire [19:0] ex_reg_rs_bypass_1_pad;
  wire [18:0] ex_reg_rs_lsb_0_shl;
  wire [19:0] ex_reg_rs_lsb_0_pad;
  wire [18:0] ex_reg_rs_lsb_1_shl;
  wire [19:0] ex_reg_rs_lsb_1_pad;
  wire [19:0] Rocket_xor32;
  wire [19:0] Rocket_xor15;
  wire [19:0] Rocket_xor34;
  wire [19:0] Rocket_xor16;
  wire [19:0] Rocket_xor7;
  wire [19:0] Rocket_xor36;
  wire [19:0] Rocket_xor17;
  wire [19:0] Rocket_xor37;
  wire [19:0] Rocket_xor38;
  wire [19:0] Rocket_xor18;
  wire [19:0] Rocket_xor8;
  wire [19:0] Rocket_xor3;
  wire [19:0] Rocket_xor40;
  wire [19:0] Rocket_xor19;
  wire [19:0] Rocket_xor42;
  wire [19:0] Rocket_xor20;
  wire [19:0] Rocket_xor9;
  wire [19:0] Rocket_xor44;
  wire [19:0] Rocket_xor21;
  wire [19:0] Rocket_xor45;
  wire [19:0] Rocket_xor46;
  wire [19:0] Rocket_xor22;
  wire [19:0] Rocket_xor10;
  wire [19:0] Rocket_xor4;
  wire [19:0] Rocket_xor1;
  wire [19:0] Rocket_xor48;
  wire [19:0] Rocket_xor23;
  wire [19:0] Rocket_xor50;
  wire [19:0] Rocket_xor24;
  wire [19:0] Rocket_xor11;
  wire [19:0] Rocket_xor52;
  wire [19:0] Rocket_xor25;
  wire [19:0] Rocket_xor53;
  wire [19:0] Rocket_xor54;
  wire [19:0] Rocket_xor26;
  wire [19:0] Rocket_xor12;
  wire [19:0] Rocket_xor5;
  wire [19:0] Rocket_xor56;
  wire [19:0] Rocket_xor27;
  wire [19:0] Rocket_xor57;
  wire [19:0] Rocket_xor58;
  wire [19:0] Rocket_xor28;
  wire [19:0] Rocket_xor13;
  wire [19:0] Rocket_xor60;
  wire [19:0] Rocket_xor29;
  wire [19:0] Rocket_xor61;
  wire [19:0] Rocket_xor62;
  wire [19:0] Rocket_xor30;
  wire [19:0] Rocket_xor14;
  wire [19:0] Rocket_xor6;
  wire [19:0] Rocket_xor2;
  wire [19:0] Rocket_xor0;
  wire [29:0] csr_sum;
  wire [29:0] div_sum;
  wire [29:0] ibuf_sum;
  wire [29:0] alu_sum;
  wire [29:0] bpu_sum;
  wire  alu_metaAssert_wire;
  wire  div_metaAssert_wire;
  wire  bpu_metaAssert_wire;
  wire  ibuf_metaAssert_wire;
  wire  csr_metaAssert_wire;
  wire  Rocket_or1;
  wire  Rocket_or6;
  wire  Rocket_or2;
  wire  Rocket_or0;
  reg  Rocket_metaAssert;
  reg [31:0] _RAND_93;
  IBuf ibuf ( // @[RocketCore.scala 236:20]
    .clock(ibuf_clock),
    .reset(ibuf_reset),
    .io_imem_ready(ibuf_io_imem_ready),
    .io_imem_valid(ibuf_io_imem_valid),
    .io_imem_bits_btb_taken(ibuf_io_imem_bits_btb_taken),
    .io_imem_bits_btb_bridx(ibuf_io_imem_bits_btb_bridx),
    .io_imem_bits_btb_entry(ibuf_io_imem_bits_btb_entry),
    .io_imem_bits_btb_bht_history(ibuf_io_imem_bits_btb_bht_history),
    .io_imem_bits_pc(ibuf_io_imem_bits_pc),
    .io_imem_bits_data(ibuf_io_imem_bits_data),
    .io_imem_bits_xcpt_pf_inst(ibuf_io_imem_bits_xcpt_pf_inst),
    .io_imem_bits_xcpt_ae_inst(ibuf_io_imem_bits_xcpt_ae_inst),
    .io_imem_bits_replay(ibuf_io_imem_bits_replay),
    .io_kill(ibuf_io_kill),
    .io_pc(ibuf_io_pc),
    .io_btb_resp_entry(ibuf_io_btb_resp_entry),
    .io_btb_resp_bht_history(ibuf_io_btb_resp_bht_history),
    .io_inst_0_ready(ibuf_io_inst_0_ready),
    .io_inst_0_valid(ibuf_io_inst_0_valid),
    .io_inst_0_bits_xcpt0_pf_inst(ibuf_io_inst_0_bits_xcpt0_pf_inst),
    .io_inst_0_bits_xcpt0_ae_inst(ibuf_io_inst_0_bits_xcpt0_ae_inst),
    .io_inst_0_bits_xcpt1_pf_inst(ibuf_io_inst_0_bits_xcpt1_pf_inst),
    .io_inst_0_bits_xcpt1_ae_inst(ibuf_io_inst_0_bits_xcpt1_ae_inst),
    .io_inst_0_bits_replay(ibuf_io_inst_0_bits_replay),
    .io_inst_0_bits_rvc(ibuf_io_inst_0_bits_rvc),
    .io_inst_0_bits_inst_bits(ibuf_io_inst_0_bits_inst_bits),
    .io_inst_0_bits_inst_rd(ibuf_io_inst_0_bits_inst_rd),
    .io_inst_0_bits_inst_rs1(ibuf_io_inst_0_bits_inst_rs1),
    .io_inst_0_bits_inst_rs2(ibuf_io_inst_0_bits_inst_rs2),
    .io_inst_0_bits_inst_rs3(ibuf_io_inst_0_bits_inst_rs3),
    .io_inst_0_bits_raw(ibuf_io_inst_0_bits_raw),
    .io_covSum(ibuf_io_covSum),
    .metaAssert(ibuf_metaAssert),
    .metaReset(ibuf_metaReset)
  );
  CSRFile csr ( // @[RocketCore.scala 257:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_ungated_clock(csr_io_ungated_clock),
    .io_interrupts_debug(csr_io_interrupts_debug),
    .io_interrupts_mtip(csr_io_interrupts_mtip),
    .io_interrupts_msip(csr_io_interrupts_msip),
    .io_interrupts_meip(csr_io_interrupts_meip),
    .io_interrupts_seip(csr_io_interrupts_seip),
    .io_hartid(csr_io_hartid),
    .io_rw_addr(csr_io_rw_addr),
    .io_rw_cmd(csr_io_rw_cmd),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_wdata(csr_io_rw_wdata),
    .io_pcode_req_valid(csr_io_pcode_req_valid),
    .io_pcode_req_bits_id(csr_io_pcode_req_bits_id),
    .io_pcode_req_bits_value_base(csr_io_pcode_req_bits_value_base),
    .io_pcode_req_bits_value_mask(csr_io_pcode_req_bits_value_mask),
    .io_pcode_req_bits_value_valid(csr_io_pcode_req_bits_value_valid),
    .io_pcode_req_bits_value_locked(csr_io_pcode_req_bits_value_locked),
    .io_vpoffset_req_bits_value(csr_io_vpoffset_req_bits_value),
    .io_decode_0_csr(csr_io_decode_0_csr),
    .io_decode_0_fp_illegal(csr_io_decode_0_fp_illegal),
    .io_decode_0_fp_csr(csr_io_decode_0_fp_csr),
    .io_decode_0_read_illegal(csr_io_decode_0_read_illegal),
    .io_decode_0_write_illegal(csr_io_decode_0_write_illegal),
    .io_decode_0_write_flush(csr_io_decode_0_write_flush),
    .io_decode_0_system_illegal(csr_io_decode_0_system_illegal),
    .io_csr_stall(csr_io_csr_stall),
    .io_eret(csr_io_eret),
    .io_singleStep(csr_io_singleStep),
    .io_status_debug(csr_io_status_debug),
    .io_status_isa(csr_io_status_isa),
    .io_status_dprv(csr_io_status_dprv),
    .io_status_prv(csr_io_status_prv),
    .io_status_sd(csr_io_status_sd),
    .io_status_zero2(csr_io_status_zero2),
    .io_status_sxl(csr_io_status_sxl),
    .io_status_uxl(csr_io_status_uxl),
    .io_status_sd_rv32(csr_io_status_sd_rv32),
    .io_status_zero1(csr_io_status_zero1),
    .io_status_tsr(csr_io_status_tsr),
    .io_status_tw(csr_io_status_tw),
    .io_status_tvm(csr_io_status_tvm),
    .io_status_mxr(csr_io_status_mxr),
    .io_status_sum(csr_io_status_sum),
    .io_status_mprv(csr_io_status_mprv),
    .io_status_xs(csr_io_status_xs),
    .io_status_fs(csr_io_status_fs),
    .io_status_mpp(csr_io_status_mpp),
    .io_status_hpp(csr_io_status_hpp),
    .io_status_spp(csr_io_status_spp),
    .io_status_mpie(csr_io_status_mpie),
    .io_status_hpie(csr_io_status_hpie),
    .io_status_spie(csr_io_status_spie),
    .io_status_upie(csr_io_status_upie),
    .io_status_mie(csr_io_status_mie),
    .io_status_hie(csr_io_status_hie),
    .io_status_sie(csr_io_status_sie),
    .io_status_uie(csr_io_status_uie),
    .io_ptbr_mode(csr_io_ptbr_mode),
    .io_ptbr_ppn(csr_io_ptbr_ppn),
    .io_evec(csr_io_evec),
    .io_exception(csr_io_exception),
    .io_retire(csr_io_retire),
    .io_cause(csr_io_cause),
    .io_pc(csr_io_pc),
    .io_tval(csr_io_tval),
    .io_fcsr_rm(csr_io_fcsr_rm),
    .io_fcsr_flags_valid(csr_io_fcsr_flags_valid),
    .io_fcsr_flags_bits(csr_io_fcsr_flags_bits),
    .io_interrupt(csr_io_interrupt),
    .io_interrupt_cause(csr_io_interrupt_cause),
    .io_bp_0_control_action(csr_io_bp_0_control_action),
    .io_bp_0_control_tmatch(csr_io_bp_0_control_tmatch),
    .io_bp_0_control_m(csr_io_bp_0_control_m),
    .io_bp_0_control_s(csr_io_bp_0_control_s),
    .io_bp_0_control_u(csr_io_bp_0_control_u),
    .io_bp_0_control_x(csr_io_bp_0_control_x),
    .io_bp_0_control_w(csr_io_bp_0_control_w),
    .io_bp_0_control_r(csr_io_bp_0_control_r),
    .io_bp_0_address(csr_io_bp_0_address),
    .io_pmp_0_cfg_l(csr_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(csr_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(csr_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(csr_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(csr_io_pmp_0_cfg_r),
    .io_pmp_0_addr(csr_io_pmp_0_addr),
    .io_pmp_0_mask(csr_io_pmp_0_mask),
    .io_pmp_1_cfg_l(csr_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(csr_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(csr_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(csr_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(csr_io_pmp_1_cfg_r),
    .io_pmp_1_addr(csr_io_pmp_1_addr),
    .io_pmp_1_mask(csr_io_pmp_1_mask),
    .io_pmp_2_cfg_l(csr_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(csr_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(csr_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(csr_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(csr_io_pmp_2_cfg_r),
    .io_pmp_2_addr(csr_io_pmp_2_addr),
    .io_pmp_2_mask(csr_io_pmp_2_mask),
    .io_pmp_3_cfg_l(csr_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(csr_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(csr_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(csr_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(csr_io_pmp_3_cfg_r),
    .io_pmp_3_addr(csr_io_pmp_3_addr),
    .io_pmp_3_mask(csr_io_pmp_3_mask),
    .io_pmp_4_cfg_l(csr_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(csr_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(csr_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(csr_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(csr_io_pmp_4_cfg_r),
    .io_pmp_4_addr(csr_io_pmp_4_addr),
    .io_pmp_4_mask(csr_io_pmp_4_mask),
    .io_pmp_5_cfg_l(csr_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(csr_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(csr_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(csr_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(csr_io_pmp_5_cfg_r),
    .io_pmp_5_addr(csr_io_pmp_5_addr),
    .io_pmp_5_mask(csr_io_pmp_5_mask),
    .io_pmp_6_cfg_l(csr_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(csr_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(csr_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(csr_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(csr_io_pmp_6_cfg_r),
    .io_pmp_6_addr(csr_io_pmp_6_addr),
    .io_pmp_6_mask(csr_io_pmp_6_mask),
    .io_pmp_7_cfg_l(csr_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(csr_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(csr_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(csr_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(csr_io_pmp_7_cfg_r),
    .io_pmp_7_addr(csr_io_pmp_7_addr),
    .io_pmp_7_mask(csr_io_pmp_7_mask),
    .io_covSum(csr_io_covSum),
    .metaAssert(csr_metaAssert),
    .metaReset(csr_metaReset)
  );
  BreakpointUnit bpu ( // @[RocketCore.scala 302:19]
    .io_status_debug(bpu_io_status_debug),
    .io_status_prv(bpu_io_status_prv),
    .io_bp_0_control_action(bpu_io_bp_0_control_action),
    .io_bp_0_control_tmatch(bpu_io_bp_0_control_tmatch),
    .io_bp_0_control_m(bpu_io_bp_0_control_m),
    .io_bp_0_control_s(bpu_io_bp_0_control_s),
    .io_bp_0_control_u(bpu_io_bp_0_control_u),
    .io_bp_0_control_x(bpu_io_bp_0_control_x),
    .io_bp_0_control_w(bpu_io_bp_0_control_w),
    .io_bp_0_control_r(bpu_io_bp_0_control_r),
    .io_bp_0_address(bpu_io_bp_0_address),
    .io_pc(bpu_io_pc),
    .io_ea(bpu_io_ea),
    .io_xcpt_if(bpu_io_xcpt_if),
    .io_xcpt_ld(bpu_io_xcpt_ld),
    .io_xcpt_st(bpu_io_xcpt_st),
    .io_debug_if(bpu_io_debug_if),
    .io_debug_ld(bpu_io_debug_ld),
    .io_debug_st(bpu_io_debug_st),
    .io_covSum(bpu_io_covSum),
    .metaAssert(bpu_metaAssert)
  );
  ALU alu ( // @[RocketCore.scala 361:19]
    .io_dw(alu_io_dw),
    .io_fn(alu_io_fn),
    .io_in2(alu_io_in2),
    .io_in1(alu_io_in1),
    .io_out(alu_io_out),
    .io_adder_out(alu_io_adder_out),
    .io_cmp_out(alu_io_cmp_out),
    .io_covSum(alu_io_covSum),
    .metaAssert(alu_metaAssert)
  );
  MulDiv div ( // @[RocketCore.scala 376:19]
    .clock(div_clock),
    .reset(div_reset),
    .io_req_ready(div_io_req_ready),
    .io_req_valid(div_io_req_valid),
    .io_req_bits_fn(div_io_req_bits_fn),
    .io_req_bits_dw(div_io_req_bits_dw),
    .io_req_bits_in1(div_io_req_bits_in1),
    .io_req_bits_in2(div_io_req_bits_in2),
    .io_req_bits_tag(div_io_req_bits_tag),
    .io_kill(div_io_kill),
    .io_resp_ready(div_io_resp_ready),
    .io_resp_valid(div_io_resp_valid),
    .io_resp_bits_data(div_io_resp_bits_data),
    .io_resp_bits_tag(div_io_resp_bits_tag),
    .io_covSum(div_io_covSum),
    .metaAssert(div_metaAssert),
    .metaReset(div_metaReset)
  );
  assign _T_760__T_767_addr = ~_T_765;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_760__T_767_data = _T_760[_T_760__T_767_addr]; // @[RocketCore.scala 932:23]
  `else
  assign _T_760__T_767_data = _T_760__T_767_addr >= 5'h1f ? _RAND_1[63:0] : _T_760[_T_760__T_767_addr]; // @[RocketCore.scala 932:23]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_760__T_775_addr = ~_T_773;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_760__T_775_data = _T_760[_T_760__T_775_addr]; // @[RocketCore.scala 932:23]
  `else
  assign _T_760__T_775_data = _T_760__T_775_addr >= 5'h1f ? _RAND_2[63:0] : _T_760[_T_760__T_775_addr]; // @[RocketCore.scala 932:23]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_760__T_1499_data = _T_1490 ? io_dmem_resp_bits_data : _T_1495;
  assign _T_760__T_1499_addr = ~rf_waddr;
  assign _T_760__T_1499_mask = 1'h1;
  assign _T_760__T_1499_en = rf_wen & _T_1496;
  assign replay_wb_common = io_dmem_s2_nack | wb_reg_replay; // @[RocketCore.scala 585:42]
  assign _T_1437 = wb_reg_valid & wb_ctrl_mem; // @[RocketCore.scala 564:19]
  assign _T_1438 = _T_1437 & io_dmem_s2_xcpt_ma_st; // @[RocketCore.scala 564:34]
  assign _T_1449 = wb_reg_xcpt | _T_1438; // @[RocketCore.scala 892:26]
  assign _T_1440 = _T_1437 & io_dmem_s2_xcpt_ma_ld; // @[RocketCore.scala 565:34]
  assign _T_1450 = _T_1449 | _T_1440; // @[RocketCore.scala 892:26]
  assign _T_1442 = _T_1437 & io_dmem_s2_xcpt_pf_st; // @[RocketCore.scala 566:34]
  assign _T_1451 = _T_1450 | _T_1442; // @[RocketCore.scala 892:26]
  assign _T_1444 = _T_1437 & io_dmem_s2_xcpt_pf_ld; // @[RocketCore.scala 567:34]
  assign _T_1452 = _T_1451 | _T_1444; // @[RocketCore.scala 892:26]
  assign _T_1446 = _T_1437 & io_dmem_s2_xcpt_ae_st; // @[RocketCore.scala 568:34]
  assign _T_1453 = _T_1452 | _T_1446; // @[RocketCore.scala 892:26]
  assign _T_1448 = _T_1437 & io_dmem_s2_xcpt_ae_ld; // @[RocketCore.scala 569:34]
  assign wb_xcpt = _T_1453 | _T_1448; // @[RocketCore.scala 892:26]
  assign _T_1475 = replay_wb_common | wb_xcpt; // @[RocketCore.scala 588:27]
  assign _T_1476 = _T_1475 | csr_io_eret; // @[RocketCore.scala 588:38]
  assign take_pc_wb = _T_1476 | wb_reg_flush_pipe; // @[RocketCore.scala 588:53]
  assign _T_1109 = ex_reg_valid | ex_reg_replay; // @[RocketCore.scala 447:34]
  assign ex_pc_valid = _T_1109 | ex_reg_xcpt_interrupt; // @[RocketCore.scala 447:51]
  assign _T_1282 = mem_ctrl_jalr | mem_reg_sfence; // @[RocketCore.scala 470:36]
  assign a = mem_reg_wdata[63:39]; // @[RocketCore.scala 906:23]
  assign _T_1284 = $signed(a) == 25'sh0; // @[RocketCore.scala 907:21]
  assign _T_1285 = $signed(a) == -25'sh1; // @[RocketCore.scala 907:34]
  assign _T_1286 = _T_1284 | _T_1285; // @[RocketCore.scala 907:29]
  assign msb = _T_1286 ? mem_reg_wdata[39] : ~mem_reg_wdata[38]; // @[RocketCore.scala 907:18]
  assign _T_1292 = {msb,mem_reg_wdata[38:0]}; // @[RocketCore.scala 470:106]
  assign _T_1152 = mem_ctrl_branch & mem_br_taken; // @[RocketCore.scala 467:25]
  assign _T_1155 = mem_reg_inst[31]; // @[RocketCore.scala 954:53]
  assign _T_1210 = mem_reg_inst[31]; // @[Cat.scala 30:58]
  assign _T_1209 = {11{_T_1155}}; // @[Cat.scala 30:58]
  assign _T_1207 = {8{_T_1155}}; // @[Cat.scala 30:58]
  assign _T_1206 = mem_reg_inst[7]; // @[Cat.scala 30:58]
  assign _T_1214 = {_T_1210,_T_1209,_T_1207,_T_1206,mem_reg_inst[30:25],mem_reg_inst[11:8],1'h0}; // @[RocketCore.scala 968:53]
  assign _T_1269 = mem_reg_inst[19:12]; // @[Cat.scala 30:58]
  assign _T_1268 = mem_reg_inst[20]; // @[Cat.scala 30:58]
  assign _T_1276 = {_T_1210,_T_1209,_T_1269,_T_1268,mem_reg_inst[30:25],mem_reg_inst[24:21],1'h0}; // @[RocketCore.scala 968:53]
  assign _T_1277 = mem_reg_rvc ? $signed(4'sh2) : $signed(4'sh4); // @[RocketCore.scala 469:8]
  assign _T_1278 = mem_ctrl_jal ? $signed(_T_1276) : $signed({{28{_T_1277[3]}},_T_1277}); // @[RocketCore.scala 468:8]
  assign _T_1279 = _T_1152 ? $signed(_T_1214) : $signed(_T_1278); // @[RocketCore.scala 467:8]
  assign _GEN_235 = {{8{_T_1279[31]}},_T_1279}; // @[RocketCore.scala 466:41]
  assign mem_br_target = $signed(mem_reg_pc) + $signed(_GEN_235); // @[RocketCore.scala 466:41]
  assign _T_1293 = _T_1282 ? $signed(_T_1292) : $signed(mem_br_target); // @[RocketCore.scala 470:21]
  assign mem_npc = $signed(_T_1293) & -40'sh2; // @[RocketCore.scala 470:141]
  assign _T_1296 = mem_npc != ex_reg_pc; // @[RocketCore.scala 472:30]
  assign _T_1297 = ibuf_io_inst_0_valid | ibuf_io_imem_valid; // @[RocketCore.scala 473:31]
  assign _T_1298 = mem_npc != ibuf_io_pc; // @[RocketCore.scala 473:62]
  assign _T_1299 = _T_1297 ? _T_1298 : 1'h1; // @[RocketCore.scala 473:8]
  assign mem_wrong_npc = ex_pc_valid ? _T_1296 : _T_1299; // @[RocketCore.scala 472:8]
  assign _T_1315 = mem_wrong_npc | mem_reg_sfence; // @[RocketCore.scala 480:54]
  assign take_pc_mem = mem_reg_valid & _T_1315; // @[RocketCore.scala 480:32]
  assign take_pc_mem_wb = take_pc_wb | take_pc_mem; // @[RocketCore.scala 232:35]
  assign _T_309 = ibuf_io_inst_0_bits_inst_bits & 32'h207f; // @[Decode.scala 14:65]
  assign _T_310 = _T_309 == 32'h3; // @[Decode.scala 14:121]
  assign _T_311 = ibuf_io_inst_0_bits_inst_bits & 32'h106f; // @[Decode.scala 14:65]
  assign _T_312 = _T_311 == 32'h3; // @[Decode.scala 14:121]
  assign _T_313 = ibuf_io_inst_0_bits_inst_bits & 32'h607f; // @[Decode.scala 14:65]
  assign _T_314 = _T_313 == 32'hf; // @[Decode.scala 14:121]
  assign _T_315 = ibuf_io_inst_0_bits_inst_bits & 32'h7077; // @[Decode.scala 14:65]
  assign _T_316 = _T_315 == 32'h13; // @[Decode.scala 14:121]
  assign _T_317 = ibuf_io_inst_0_bits_inst_bits & 32'h5f; // @[Decode.scala 14:65]
  assign _T_318 = _T_317 == 32'h17; // @[Decode.scala 14:121]
  assign _T_319 = ibuf_io_inst_0_bits_inst_bits & 32'hfc00007f; // @[Decode.scala 14:65]
  assign _T_320 = _T_319 == 32'h33; // @[Decode.scala 14:121]
  assign _T_321 = ibuf_io_inst_0_bits_inst_bits & 32'hbe007077; // @[Decode.scala 14:65]
  assign _T_322 = _T_321 == 32'h33; // @[Decode.scala 14:121]
  assign _T_323 = ibuf_io_inst_0_bits_inst_bits & 32'h4000073; // @[Decode.scala 14:65]
  assign _T_324 = _T_323 == 32'h43; // @[Decode.scala 14:121]
  assign _T_325 = ibuf_io_inst_0_bits_inst_bits & 32'he400007f; // @[Decode.scala 14:65]
  assign _T_326 = _T_325 == 32'h53; // @[Decode.scala 14:121]
  assign _T_327 = ibuf_io_inst_0_bits_inst_bits & 32'h707b; // @[Decode.scala 14:65]
  assign _T_328 = _T_327 == 32'h63; // @[Decode.scala 14:121]
  assign _T_329 = ibuf_io_inst_0_bits_inst_bits & 32'h7f; // @[Decode.scala 14:65]
  assign _T_330 = _T_329 == 32'h6f; // @[Decode.scala 14:121]
  assign _T_331 = ibuf_io_inst_0_bits_inst_bits & 32'hffefffff; // @[Decode.scala 14:65]
  assign _T_332 = _T_331 == 32'h73; // @[Decode.scala 14:121]
  assign _T_333 = ibuf_io_inst_0_bits_inst_bits & 32'hfc00305f; // @[Decode.scala 14:65]
  assign _T_334 = _T_333 == 32'h1013; // @[Decode.scala 14:121]
  assign _T_335 = ibuf_io_inst_0_bits_inst_bits & 32'hfe00305f; // @[Decode.scala 14:65]
  assign _T_336 = _T_335 == 32'h101b; // @[Decode.scala 14:121]
  assign _T_337 = ibuf_io_inst_0_bits_inst_bits & 32'h605b; // @[Decode.scala 14:65]
  assign _T_338 = _T_337 == 32'h2003; // @[Decode.scala 14:121]
  assign _T_340 = _T_309 == 32'h2013; // @[Decode.scala 14:121]
  assign _T_341 = ibuf_io_inst_0_bits_inst_bits & 32'h1800607f; // @[Decode.scala 14:65]
  assign _T_342 = _T_341 == 32'h202f; // @[Decode.scala 14:121]
  assign _T_344 = _T_309 == 32'h2073; // @[Decode.scala 14:121]
  assign _T_345 = ibuf_io_inst_0_bits_inst_bits & 32'hbc00707f; // @[Decode.scala 14:65]
  assign _T_346 = _T_345 == 32'h5013; // @[Decode.scala 14:121]
  assign _T_347 = ibuf_io_inst_0_bits_inst_bits & 32'hbe00705f; // @[Decode.scala 14:65]
  assign _T_348 = _T_347 == 32'h501b; // @[Decode.scala 14:121]
  assign _T_350 = _T_321 == 32'h5033; // @[Decode.scala 14:121]
  assign _T_351 = ibuf_io_inst_0_bits_inst_bits & 32'hfe004077; // @[Decode.scala 14:65]
  assign _T_352 = _T_351 == 32'h2004033; // @[Decode.scala 14:121]
  assign _T_353 = ibuf_io_inst_0_bits_inst_bits & 32'he800607f; // @[Decode.scala 14:65]
  assign _T_354 = _T_353 == 32'h800202f; // @[Decode.scala 14:121]
  assign _T_355 = ibuf_io_inst_0_bits_inst_bits & 32'hf9f0607f; // @[Decode.scala 14:65]
  assign _T_356 = _T_355 == 32'h1000202f; // @[Decode.scala 14:121]
  assign _T_357 = ibuf_io_inst_0_bits_inst_bits & 32'hdfffffff; // @[Decode.scala 14:65]
  assign _T_358 = _T_357 == 32'h10200073; // @[Decode.scala 14:121]
  assign _T_359 = ibuf_io_inst_0_bits_inst_bits == 32'h10500073; // @[Decode.scala 14:121]
  assign _T_360 = ibuf_io_inst_0_bits_inst_bits & 32'hfe007fff; // @[Decode.scala 14:65]
  assign _T_361 = _T_360 == 32'h12000073; // @[Decode.scala 14:121]
  assign _T_362 = ibuf_io_inst_0_bits_inst_bits & 32'hf400607f; // @[Decode.scala 14:65]
  assign _T_363 = _T_362 == 32'h20000053; // @[Decode.scala 14:121]
  assign _T_364 = ibuf_io_inst_0_bits_inst_bits & 32'h7c00607f; // @[Decode.scala 14:65]
  assign _T_365 = _T_364 == 32'h20000053; // @[Decode.scala 14:121]
  assign _T_366 = ibuf_io_inst_0_bits_inst_bits & 32'h7c00507f; // @[Decode.scala 14:65]
  assign _T_367 = _T_366 == 32'h20000053; // @[Decode.scala 14:121]
  assign _T_368 = ibuf_io_inst_0_bits_inst_bits & 32'h7ff0007f; // @[Decode.scala 14:65]
  assign _T_369 = _T_368 == 32'h40100053; // @[Decode.scala 14:121]
  assign _T_371 = _T_368 == 32'h42000053; // @[Decode.scala 14:121]
  assign _T_372 = ibuf_io_inst_0_bits_inst_bits & 32'hfdf0007f; // @[Decode.scala 14:65]
  assign _T_373 = _T_372 == 32'h58000053; // @[Decode.scala 14:121]
  assign _T_374 = ibuf_io_inst_0_bits_inst_bits == 32'h7b200073; // @[Decode.scala 14:121]
  assign _T_375 = ibuf_io_inst_0_bits_inst_bits & 32'hedc0007f; // @[Decode.scala 14:65]
  assign _T_376 = _T_375 == 32'hc0000053; // @[Decode.scala 14:121]
  assign _T_377 = ibuf_io_inst_0_bits_inst_bits & 32'hfdf0607f; // @[Decode.scala 14:65]
  assign _T_378 = _T_377 == 32'he0000053; // @[Decode.scala 14:121]
  assign _T_379 = ibuf_io_inst_0_bits_inst_bits & 32'hedf0707f; // @[Decode.scala 14:65]
  assign _T_380 = _T_379 == 32'he0000053; // @[Decode.scala 14:121]
  assign _T_381 = ibuf_io_inst_0_bits_inst_bits & 32'h306f; // @[Decode.scala 14:65]
  assign _T_382 = _T_381 == 32'h1063; // @[Decode.scala 14:121]
  assign _T_383 = ibuf_io_inst_0_bits_inst_bits & 32'h407f; // @[Decode.scala 14:65]
  assign _T_384 = _T_383 == 32'h4063; // @[Decode.scala 14:121]
  assign _T_385 = ibuf_io_inst_0_bits_inst_bits & 32'hfc007077; // @[Decode.scala 14:65]
  assign _T_386 = _T_385 == 32'h33; // @[Decode.scala 14:121]
  assign _T_387 = ibuf_io_inst_0_bits_inst_bits & 32'h405f; // @[Decode.scala 14:65]
  assign _T_388 = _T_387 == 32'h3; // @[Decode.scala 14:121]
  assign _T_390 = _T_310 | _T_312; // @[Decode.scala 15:30]
  assign _T_391 = _T_390 | _T_314; // @[Decode.scala 15:30]
  assign _T_392 = _T_391 | _T_316; // @[Decode.scala 15:30]
  assign _T_393 = _T_392 | _T_318; // @[Decode.scala 15:30]
  assign _T_394 = _T_393 | _T_320; // @[Decode.scala 15:30]
  assign _T_395 = _T_394 | _T_322; // @[Decode.scala 15:30]
  assign _T_396 = _T_395 | _T_324; // @[Decode.scala 15:30]
  assign _T_397 = _T_396 | _T_326; // @[Decode.scala 15:30]
  assign _T_398 = _T_397 | _T_328; // @[Decode.scala 15:30]
  assign _T_399 = _T_398 | _T_330; // @[Decode.scala 15:30]
  assign _T_400 = _T_399 | _T_332; // @[Decode.scala 15:30]
  assign _T_401 = _T_400 | _T_334; // @[Decode.scala 15:30]
  assign _T_402 = _T_401 | _T_336; // @[Decode.scala 15:30]
  assign _T_403 = _T_402 | _T_338; // @[Decode.scala 15:30]
  assign _T_404 = _T_403 | _T_340; // @[Decode.scala 15:30]
  assign _T_405 = _T_404 | _T_342; // @[Decode.scala 15:30]
  assign _T_406 = _T_405 | _T_344; // @[Decode.scala 15:30]
  assign _T_407 = _T_406 | _T_346; // @[Decode.scala 15:30]
  assign _T_408 = _T_407 | _T_348; // @[Decode.scala 15:30]
  assign _T_409 = _T_408 | _T_350; // @[Decode.scala 15:30]
  assign _T_410 = _T_409 | _T_352; // @[Decode.scala 15:30]
  assign _T_411 = _T_410 | _T_354; // @[Decode.scala 15:30]
  assign _T_412 = _T_411 | _T_356; // @[Decode.scala 15:30]
  assign _T_413 = _T_412 | _T_358; // @[Decode.scala 15:30]
  assign _T_414 = _T_413 | _T_359; // @[Decode.scala 15:30]
  assign _T_415 = _T_414 | _T_361; // @[Decode.scala 15:30]
  assign _T_416 = _T_415 | _T_363; // @[Decode.scala 15:30]
  assign _T_417 = _T_416 | _T_365; // @[Decode.scala 15:30]
  assign _T_418 = _T_417 | _T_367; // @[Decode.scala 15:30]
  assign _T_419 = _T_418 | _T_369; // @[Decode.scala 15:30]
  assign _T_420 = _T_419 | _T_371; // @[Decode.scala 15:30]
  assign _T_421 = _T_420 | _T_373; // @[Decode.scala 15:30]
  assign _T_422 = _T_421 | _T_374; // @[Decode.scala 15:30]
  assign _T_423 = _T_422 | _T_376; // @[Decode.scala 15:30]
  assign _T_424 = _T_423 | _T_378; // @[Decode.scala 15:30]
  assign _T_425 = _T_424 | _T_380; // @[Decode.scala 15:30]
  assign _T_426 = _T_425 | _T_382; // @[Decode.scala 15:30]
  assign _T_427 = _T_426 | _T_384; // @[Decode.scala 15:30]
  assign _T_428 = _T_427 | _T_386; // @[Decode.scala 15:30]
  assign id_ctrl_legal = _T_428 | _T_388; // @[Decode.scala 15:30]
  assign _T_430 = ibuf_io_inst_0_bits_inst_bits & 32'h5c; // @[Decode.scala 14:65]
  assign _T_431 = _T_430 == 32'h4; // @[Decode.scala 14:121]
  assign _T_432 = ibuf_io_inst_0_bits_inst_bits & 32'h60; // @[Decode.scala 14:65]
  assign _T_433 = _T_432 == 32'h40; // @[Decode.scala 14:121]
  assign id_ctrl_fp = _T_431 | _T_433; // @[Decode.scala 15:30]
  assign _T_436 = ibuf_io_inst_0_bits_inst_bits & 32'h74; // @[Decode.scala 14:65]
  assign id_ctrl_branch = _T_436 == 32'h60; // @[Decode.scala 14:121]
  assign _T_439 = ibuf_io_inst_0_bits_inst_bits & 32'h68; // @[Decode.scala 14:65]
  assign id_ctrl_jal = _T_439 == 32'h68; // @[Decode.scala 14:121]
  assign _T_442 = ibuf_io_inst_0_bits_inst_bits & 32'h203c; // @[Decode.scala 14:65]
  assign id_ctrl_jalr = _T_442 == 32'h24; // @[Decode.scala 14:121]
  assign _T_445 = ibuf_io_inst_0_bits_inst_bits & 32'h64; // @[Decode.scala 14:65]
  assign _T_446 = _T_445 == 32'h20; // @[Decode.scala 14:121]
  assign _T_447 = ibuf_io_inst_0_bits_inst_bits & 32'h34; // @[Decode.scala 14:65]
  assign _T_448 = _T_447 == 32'h20; // @[Decode.scala 14:121]
  assign _T_449 = ibuf_io_inst_0_bits_inst_bits & 32'h2048; // @[Decode.scala 14:65]
  assign _T_450 = _T_449 == 32'h2008; // @[Decode.scala 14:121]
  assign _T_451 = ibuf_io_inst_0_bits_inst_bits & 32'h42003024; // @[Decode.scala 14:65]
  assign _T_452 = _T_451 == 32'h2000020; // @[Decode.scala 14:121]
  assign _T_454 = _T_446 | _T_448; // @[Decode.scala 15:30]
  assign _T_455 = _T_454 | _T_450; // @[Decode.scala 15:30]
  assign id_ctrl_rxs2 = _T_455 | _T_452; // @[Decode.scala 15:30]
  assign _T_457 = ibuf_io_inst_0_bits_inst_bits & 32'h44; // @[Decode.scala 14:65]
  assign _T_458 = _T_457 == 32'h0; // @[Decode.scala 14:121]
  assign _T_459 = ibuf_io_inst_0_bits_inst_bits & 32'h4024; // @[Decode.scala 14:65]
  assign _T_460 = _T_459 == 32'h20; // @[Decode.scala 14:121]
  assign _T_461 = ibuf_io_inst_0_bits_inst_bits & 32'h38; // @[Decode.scala 14:65]
  assign _T_462 = _T_461 == 32'h20; // @[Decode.scala 14:121]
  assign _T_463 = ibuf_io_inst_0_bits_inst_bits & 32'h2050; // @[Decode.scala 14:65]
  assign _T_464 = _T_463 == 32'h2000; // @[Decode.scala 14:121]
  assign _T_465 = ibuf_io_inst_0_bits_inst_bits & 32'h90000034; // @[Decode.scala 14:65]
  assign _T_466 = _T_465 == 32'h90000010; // @[Decode.scala 14:121]
  assign _T_468 = _T_458 | _T_460; // @[Decode.scala 15:30]
  assign _T_469 = _T_468 | _T_462; // @[Decode.scala 15:30]
  assign _T_470 = _T_469 | _T_464; // @[Decode.scala 15:30]
  assign id_ctrl_rxs1 = _T_470 | _T_466; // @[Decode.scala 15:30]
  assign _T_472 = ibuf_io_inst_0_bits_inst_bits & 32'h58; // @[Decode.scala 14:65]
  assign _T_473 = _T_472 == 32'h0; // @[Decode.scala 14:121]
  assign _T_474 = ibuf_io_inst_0_bits_inst_bits & 32'h20; // @[Decode.scala 14:65]
  assign _T_475 = _T_474 == 32'h0; // @[Decode.scala 14:121]
  assign _T_476 = ibuf_io_inst_0_bits_inst_bits & 32'hc; // @[Decode.scala 14:65]
  assign _T_477 = _T_476 == 32'h4; // @[Decode.scala 14:121]
  assign _T_478 = ibuf_io_inst_0_bits_inst_bits & 32'h48; // @[Decode.scala 14:65]
  assign _T_479 = _T_478 == 32'h48; // @[Decode.scala 14:121]
  assign _T_480 = ibuf_io_inst_0_bits_inst_bits & 32'h4050; // @[Decode.scala 14:65]
  assign _T_481 = _T_480 == 32'h4050; // @[Decode.scala 14:121]
  assign _T_483 = _T_473 | _T_475; // @[Decode.scala 15:30]
  assign _T_484 = _T_483 | _T_477; // @[Decode.scala 15:30]
  assign _T_485 = _T_484 | _T_479; // @[Decode.scala 15:30]
  assign _T_486 = _T_485 | _T_481; // @[Decode.scala 15:30]
  assign _T_488 = _T_478 == 32'h0; // @[Decode.scala 14:121]
  assign _T_489 = ibuf_io_inst_0_bits_inst_bits & 32'h18; // @[Decode.scala 14:65]
  assign _T_490 = _T_489 == 32'h0; // @[Decode.scala 14:121]
  assign _T_491 = ibuf_io_inst_0_bits_inst_bits & 32'h4008; // @[Decode.scala 14:65]
  assign _T_492 = _T_491 == 32'h4000; // @[Decode.scala 14:121]
  assign _T_494 = _T_488 | _T_458; // @[Decode.scala 15:30]
  assign _T_495 = _T_494 | _T_490; // @[Decode.scala 15:30]
  assign _T_496 = _T_495 | _T_492; // @[Decode.scala 15:30]
  assign id_ctrl_sel_alu2 = {_T_496,_T_486}; // @[Cat.scala 30:58]
  assign _T_498 = ibuf_io_inst_0_bits_inst_bits & 32'h4004; // @[Decode.scala 14:65]
  assign _T_499 = _T_498 == 32'h0; // @[Decode.scala 14:121]
  assign _T_500 = ibuf_io_inst_0_bits_inst_bits & 32'h50; // @[Decode.scala 14:65]
  assign _T_501 = _T_500 == 32'h0; // @[Decode.scala 14:121]
  assign _T_502 = ibuf_io_inst_0_bits_inst_bits & 32'h24; // @[Decode.scala 14:65]
  assign _T_503 = _T_502 == 32'h0; // @[Decode.scala 14:121]
  assign _T_505 = _T_499 | _T_501; // @[Decode.scala 15:30]
  assign _T_506 = _T_505 | _T_458; // @[Decode.scala 15:30]
  assign _T_507 = _T_506 | _T_503; // @[Decode.scala 15:30]
  assign _T_508 = _T_507 | _T_490; // @[Decode.scala 15:30]
  assign _T_510 = _T_447 == 32'h14; // @[Decode.scala 14:121]
  assign _T_512 = _T_510 | _T_479; // @[Decode.scala 15:30]
  assign id_ctrl_sel_alu1 = {_T_512,_T_508}; // @[Cat.scala 30:58]
  assign _T_515 = _T_489 == 32'h8; // @[Decode.scala 14:121]
  assign _T_517 = _T_457 == 32'h40; // @[Decode.scala 14:121]
  assign _T_519 = _T_515 | _T_517; // @[Decode.scala 15:30]
  assign _T_520 = ibuf_io_inst_0_bits_inst_bits & 32'h14; // @[Decode.scala 14:65]
  assign _T_521 = _T_520 == 32'h14; // @[Decode.scala 14:121]
  assign _T_523 = _T_515 | _T_521; // @[Decode.scala 15:30]
  assign _T_524 = ibuf_io_inst_0_bits_inst_bits & 32'h30; // @[Decode.scala 14:65]
  assign _T_525 = _T_524 == 32'h0; // @[Decode.scala 14:121]
  assign _T_526 = ibuf_io_inst_0_bits_inst_bits & 32'h201c; // @[Decode.scala 14:65]
  assign _T_527 = _T_526 == 32'h4; // @[Decode.scala 14:121]
  assign _T_529 = _T_520 == 32'h10; // @[Decode.scala 14:121]
  assign _T_531 = _T_525 | _T_527; // @[Decode.scala 15:30]
  assign _T_532 = _T_531 | _T_529; // @[Decode.scala 15:30]
  assign id_ctrl_sel_imm = {_T_532,_T_523,_T_519}; // @[Cat.scala 30:58]
  assign _T_535 = ibuf_io_inst_0_bits_inst_bits & 32'h10; // @[Decode.scala 14:65]
  assign _T_536 = _T_535 == 32'h0; // @[Decode.scala 14:121]
  assign _T_537 = ibuf_io_inst_0_bits_inst_bits & 32'h8; // @[Decode.scala 14:65]
  assign _T_538 = _T_537 == 32'h0; // @[Decode.scala 14:121]
  assign id_ctrl_alu_dw = _T_536 | _T_538; // @[Decode.scala 15:30]
  assign _T_541 = ibuf_io_inst_0_bits_inst_bits & 32'h3054; // @[Decode.scala 14:65]
  assign _T_542 = _T_541 == 32'h1010; // @[Decode.scala 14:121]
  assign _T_543 = ibuf_io_inst_0_bits_inst_bits & 32'h1058; // @[Decode.scala 14:65]
  assign _T_544 = _T_543 == 32'h1040; // @[Decode.scala 14:121]
  assign _T_545 = ibuf_io_inst_0_bits_inst_bits & 32'h7044; // @[Decode.scala 14:65]
  assign _T_546 = _T_545 == 32'h7000; // @[Decode.scala 14:121]
  assign _T_547 = ibuf_io_inst_0_bits_inst_bits & 32'h2001074; // @[Decode.scala 14:65]
  assign _T_548 = _T_547 == 32'h2001030; // @[Decode.scala 14:121]
  assign _T_550 = _T_542 | _T_544; // @[Decode.scala 15:30]
  assign _T_551 = _T_550 | _T_546; // @[Decode.scala 15:30]
  assign _T_552 = _T_551 | _T_548; // @[Decode.scala 15:30]
  assign _T_553 = ibuf_io_inst_0_bits_inst_bits & 32'h4054; // @[Decode.scala 14:65]
  assign _T_554 = _T_553 == 32'h40; // @[Decode.scala 14:121]
  assign _T_555 = ibuf_io_inst_0_bits_inst_bits & 32'h2058; // @[Decode.scala 14:65]
  assign _T_556 = _T_555 == 32'h2040; // @[Decode.scala 14:121]
  assign _T_558 = _T_541 == 32'h3010; // @[Decode.scala 14:121]
  assign _T_559 = ibuf_io_inst_0_bits_inst_bits & 32'h6054; // @[Decode.scala 14:65]
  assign _T_560 = _T_559 == 32'h6010; // @[Decode.scala 14:121]
  assign _T_561 = ibuf_io_inst_0_bits_inst_bits & 32'h2002074; // @[Decode.scala 14:65]
  assign _T_562 = _T_561 == 32'h2002030; // @[Decode.scala 14:121]
  assign _T_563 = ibuf_io_inst_0_bits_inst_bits & 32'h40003034; // @[Decode.scala 14:65]
  assign _T_564 = _T_563 == 32'h40000030; // @[Decode.scala 14:121]
  assign _T_565 = ibuf_io_inst_0_bits_inst_bits & 32'h40001054; // @[Decode.scala 14:65]
  assign _T_566 = _T_565 == 32'h40001010; // @[Decode.scala 14:121]
  assign _T_568 = _T_554 | _T_556; // @[Decode.scala 15:30]
  assign _T_569 = _T_568 | _T_558; // @[Decode.scala 15:30]
  assign _T_570 = _T_569 | _T_560; // @[Decode.scala 15:30]
  assign _T_571 = _T_570 | _T_562; // @[Decode.scala 15:30]
  assign _T_572 = _T_571 | _T_564; // @[Decode.scala 15:30]
  assign _T_573 = _T_572 | _T_566; // @[Decode.scala 15:30]
  assign _T_574 = ibuf_io_inst_0_bits_inst_bits & 32'h2002054; // @[Decode.scala 14:65]
  assign _T_575 = _T_574 == 32'h2010; // @[Decode.scala 14:121]
  assign _T_576 = ibuf_io_inst_0_bits_inst_bits & 32'h2034; // @[Decode.scala 14:65]
  assign _T_577 = _T_576 == 32'h2010; // @[Decode.scala 14:121]
  assign _T_578 = ibuf_io_inst_0_bits_inst_bits & 32'h40004054; // @[Decode.scala 14:65]
  assign _T_579 = _T_578 == 32'h4010; // @[Decode.scala 14:121]
  assign _T_580 = ibuf_io_inst_0_bits_inst_bits & 32'h5054; // @[Decode.scala 14:65]
  assign _T_581 = _T_580 == 32'h4010; // @[Decode.scala 14:121]
  assign _T_582 = ibuf_io_inst_0_bits_inst_bits & 32'h4058; // @[Decode.scala 14:65]
  assign _T_583 = _T_582 == 32'h4040; // @[Decode.scala 14:121]
  assign _T_585 = _T_575 | _T_577; // @[Decode.scala 15:30]
  assign _T_586 = _T_585 | _T_579; // @[Decode.scala 15:30]
  assign _T_587 = _T_586 | _T_581; // @[Decode.scala 15:30]
  assign _T_588 = _T_587 | _T_583; // @[Decode.scala 15:30]
  assign _T_589 = ibuf_io_inst_0_bits_inst_bits & 32'h2006054; // @[Decode.scala 14:65]
  assign _T_590 = _T_589 == 32'h2010; // @[Decode.scala 14:121]
  assign _T_591 = ibuf_io_inst_0_bits_inst_bits & 32'h6034; // @[Decode.scala 14:65]
  assign _T_592 = _T_591 == 32'h2010; // @[Decode.scala 14:121]
  assign _T_593 = ibuf_io_inst_0_bits_inst_bits & 32'h40003054; // @[Decode.scala 14:65]
  assign _T_594 = _T_593 == 32'h40001010; // @[Decode.scala 14:121]
  assign _T_596 = _T_590 | _T_592; // @[Decode.scala 15:30]
  assign _T_597 = _T_596 | _T_583; // @[Decode.scala 15:30]
  assign _T_598 = _T_597 | _T_564; // @[Decode.scala 15:30]
  assign _T_599 = _T_598 | _T_594; // @[Decode.scala 15:30]
  assign id_ctrl_alu_fn = {_T_599,_T_588,_T_573,_T_552}; // @[Cat.scala 30:58]
  assign _T_603 = ibuf_io_inst_0_bits_inst_bits & 32'h107f; // @[Decode.scala 14:65]
  assign _T_604 = _T_603 == 32'h3; // @[Decode.scala 14:121]
  assign _T_605 = ibuf_io_inst_0_bits_inst_bits & 32'h707f; // @[Decode.scala 14:65]
  assign _T_606 = _T_605 == 32'h100f; // @[Decode.scala 14:121]
  assign _T_608 = _T_388 | _T_310; // @[Decode.scala 15:30]
  assign _T_609 = _T_608 | _T_604; // @[Decode.scala 15:30]
  assign _T_610 = _T_609 | _T_606; // @[Decode.scala 15:30]
  assign _T_611 = _T_610 | _T_338; // @[Decode.scala 15:30]
  assign _T_612 = _T_611 | _T_342; // @[Decode.scala 15:30]
  assign _T_613 = _T_612 | _T_354; // @[Decode.scala 15:30]
  assign _T_614 = _T_613 | _T_356; // @[Decode.scala 15:30]
  assign id_ctrl_mem = _T_614 | _T_361; // @[Decode.scala 15:30]
  assign _T_616 = ibuf_io_inst_0_bits_inst_bits & 32'h2008; // @[Decode.scala 14:65]
  assign _T_617 = _T_616 == 32'h8; // @[Decode.scala 14:121]
  assign _T_619 = _T_439 == 32'h20; // @[Decode.scala 14:121]
  assign _T_620 = ibuf_io_inst_0_bits_inst_bits & 32'h18000020; // @[Decode.scala 14:65]
  assign _T_621 = _T_620 == 32'h18000020; // @[Decode.scala 14:121]
  assign _T_622 = ibuf_io_inst_0_bits_inst_bits & 32'h20000020; // @[Decode.scala 14:65]
  assign _T_623 = _T_622 == 32'h20000020; // @[Decode.scala 14:121]
  assign _T_625 = _T_617 | _T_619; // @[Decode.scala 15:30]
  assign _T_626 = _T_625 | _T_621; // @[Decode.scala 15:30]
  assign _T_627 = _T_626 | _T_623; // @[Decode.scala 15:30]
  assign _T_628 = ibuf_io_inst_0_bits_inst_bits & 32'h10002008; // @[Decode.scala 14:65]
  assign _T_629 = _T_628 == 32'h10002008; // @[Decode.scala 14:121]
  assign _T_630 = ibuf_io_inst_0_bits_inst_bits & 32'h40002008; // @[Decode.scala 14:65]
  assign _T_631 = _T_630 == 32'h40002008; // @[Decode.scala 14:121]
  assign _T_633 = _T_629 | _T_631; // @[Decode.scala 15:30]
  assign _T_634 = ibuf_io_inst_0_bits_inst_bits & 32'h40; // @[Decode.scala 14:65]
  assign _T_635 = _T_634 == 32'h40; // @[Decode.scala 14:121]
  assign _T_636 = ibuf_io_inst_0_bits_inst_bits & 32'h8000008; // @[Decode.scala 14:65]
  assign _T_637 = _T_636 == 32'h8000008; // @[Decode.scala 14:121]
  assign _T_638 = ibuf_io_inst_0_bits_inst_bits & 32'h10000008; // @[Decode.scala 14:65]
  assign _T_639 = _T_638 == 32'h10000008; // @[Decode.scala 14:121]
  assign _T_640 = ibuf_io_inst_0_bits_inst_bits & 32'h80000008; // @[Decode.scala 14:65]
  assign _T_641 = _T_640 == 32'h80000008; // @[Decode.scala 14:121]
  assign _T_643 = _T_617 | _T_635; // @[Decode.scala 15:30]
  assign _T_644 = _T_643 | _T_637; // @[Decode.scala 15:30]
  assign _T_645 = _T_644 | _T_639; // @[Decode.scala 15:30]
  assign _T_646 = _T_645 | _T_641; // @[Decode.scala 15:30]
  assign _T_647 = ibuf_io_inst_0_bits_inst_bits & 32'h18002008; // @[Decode.scala 14:65]
  assign _T_648 = _T_647 == 32'h2008; // @[Decode.scala 14:121]
  assign id_ctrl_mem_cmd = {_T_635,_T_648,_T_646,_T_633,_T_627}; // @[Cat.scala 30:58]
  assign _T_655 = ibuf_io_inst_0_bits_inst_bits & 32'h1000; // @[Decode.scala 14:65]
  assign _T_656 = _T_655 == 32'h1000; // @[Decode.scala 14:121]
  assign _T_658 = ibuf_io_inst_0_bits_inst_bits & 32'h2000; // @[Decode.scala 14:65]
  assign _T_659 = _T_658 == 32'h2000; // @[Decode.scala 14:121]
  assign _T_661 = _T_635 | _T_659; // @[Decode.scala 15:30]
  assign _T_662 = ibuf_io_inst_0_bits_inst_bits & 32'h4000; // @[Decode.scala 14:65]
  assign _T_663 = _T_662 == 32'h4000; // @[Decode.scala 14:121]
  assign id_ctrl_mem_type = {_T_663,_T_661,_T_656}; // @[Cat.scala 30:58]
  assign _T_667 = ibuf_io_inst_0_bits_inst_bits & 32'h80000060; // @[Decode.scala 14:65]
  assign _T_668 = _T_667 == 32'h40; // @[Decode.scala 14:121]
  assign _T_669 = ibuf_io_inst_0_bits_inst_bits & 32'h10000060; // @[Decode.scala 14:65]
  assign _T_671 = ibuf_io_inst_0_bits_inst_bits & 32'h70; // @[Decode.scala 14:65]
  assign id_ctrl_rfs3 = _T_671 == 32'h40; // @[Decode.scala 14:121]
  assign _T_687 = ibuf_io_inst_0_bits_inst_bits & 32'h3c; // @[Decode.scala 14:65]
  assign _T_688 = _T_687 == 32'h4; // @[Decode.scala 14:121]
  assign _T_690 = _T_669 == 32'h10000040; // @[Decode.scala 14:121]
  assign _T_692 = _T_688 | _T_668; // @[Decode.scala 15:30]
  assign _T_693 = _T_692 | id_ctrl_rfs3; // @[Decode.scala 15:30]
  assign id_ctrl_wfd = _T_693 | _T_690; // @[Decode.scala 15:30]
  assign _T_695 = ibuf_io_inst_0_bits_inst_bits & 32'h2000074; // @[Decode.scala 14:65]
  assign id_ctrl_div = _T_695 == 32'h2000030; // @[Decode.scala 14:121]
  assign _T_699 = _T_445 == 32'h0; // @[Decode.scala 14:121]
  assign _T_701 = _T_500 == 32'h10; // @[Decode.scala 14:121]
  assign _T_702 = ibuf_io_inst_0_bits_inst_bits & 32'h2024; // @[Decode.scala 14:65]
  assign _T_703 = _T_702 == 32'h24; // @[Decode.scala 14:121]
  assign _T_704 = ibuf_io_inst_0_bits_inst_bits & 32'h28; // @[Decode.scala 14:65]
  assign _T_705 = _T_704 == 32'h28; // @[Decode.scala 14:121]
  assign _T_706 = ibuf_io_inst_0_bits_inst_bits & 32'h1030; // @[Decode.scala 14:65]
  assign _T_707 = _T_706 == 32'h1030; // @[Decode.scala 14:121]
  assign _T_708 = ibuf_io_inst_0_bits_inst_bits & 32'h2030; // @[Decode.scala 14:65]
  assign _T_709 = _T_708 == 32'h2030; // @[Decode.scala 14:121]
  assign _T_710 = ibuf_io_inst_0_bits_inst_bits & 32'h90000010; // @[Decode.scala 14:65]
  assign _T_711 = _T_710 == 32'h80000010; // @[Decode.scala 14:121]
  assign _T_713 = _T_699 | _T_701; // @[Decode.scala 15:30]
  assign _T_714 = _T_713 | _T_703; // @[Decode.scala 15:30]
  assign _T_715 = _T_714 | _T_705; // @[Decode.scala 15:30]
  assign _T_716 = _T_715 | _T_707; // @[Decode.scala 15:30]
  assign _T_717 = _T_716 | _T_709; // @[Decode.scala 15:30]
  assign id_ctrl_wxd = _T_717 | _T_711; // @[Decode.scala 15:30]
  assign _T_719 = ibuf_io_inst_0_bits_inst_bits & 32'h1070; // @[Decode.scala 14:65]
  assign _T_720 = _T_719 == 32'h1070; // @[Decode.scala 14:121]
  assign _T_722 = ibuf_io_inst_0_bits_inst_bits & 32'h2070; // @[Decode.scala 14:65]
  assign _T_723 = _T_722 == 32'h2070; // @[Decode.scala 14:121]
  assign _T_725 = ibuf_io_inst_0_bits_inst_bits & 32'h10000070; // @[Decode.scala 14:65]
  assign _T_726 = _T_725 == 32'h70; // @[Decode.scala 14:121]
  assign _T_727 = ibuf_io_inst_0_bits_inst_bits & 32'h12000034; // @[Decode.scala 14:65]
  assign _T_728 = _T_727 == 32'h10000030; // @[Decode.scala 14:121]
  assign _T_729 = ibuf_io_inst_0_bits_inst_bits & 32'he0000050; // @[Decode.scala 14:65]
  assign _T_730 = _T_729 == 32'h60000050; // @[Decode.scala 14:121]
  assign _T_732 = _T_726 | _T_720; // @[Decode.scala 15:30]
  assign _T_733 = _T_732 | _T_723; // @[Decode.scala 15:30]
  assign _T_734 = _T_733 | _T_728; // @[Decode.scala 15:30]
  assign _T_735 = _T_734 | _T_730; // @[Decode.scala 15:30]
  assign id_ctrl_csr = {_T_735,_T_723,_T_720}; // @[Cat.scala 30:58]
  assign _T_738 = ibuf_io_inst_0_bits_inst_bits & 32'h3058; // @[Decode.scala 14:65]
  assign id_ctrl_fence_i = _T_738 == 32'h1008; // @[Decode.scala 14:121]
  assign id_ctrl_fence = _T_738 == 32'h8; // @[Decode.scala 14:121]
  assign _T_744 = ibuf_io_inst_0_bits_inst_bits & 32'h6048; // @[Decode.scala 14:65]
  assign id_ctrl_amo = _T_744 == 32'h2008; // @[Decode.scala 14:121]
  assign _T_747 = ibuf_io_inst_0_bits_inst_bits & 32'h105c; // @[Decode.scala 14:65]
  assign _T_748 = _T_747 == 32'h1004; // @[Decode.scala 14:121]
  assign _T_749 = ibuf_io_inst_0_bits_inst_bits & 32'h2000060; // @[Decode.scala 14:65]
  assign _T_750 = _T_749 == 32'h2000040; // @[Decode.scala 14:121]
  assign _T_751 = ibuf_io_inst_0_bits_inst_bits & 32'hd0000070; // @[Decode.scala 14:65]
  assign _T_752 = _T_751 == 32'h40000050; // @[Decode.scala 14:121]
  assign _T_754 = _T_748 | _T_750; // @[Decode.scala 15:30]
  assign id_ctrl_dp = _T_754 | _T_752; // @[Decode.scala 15:30]
  assign _T_763 = ibuf_io_inst_0_bits_inst_rs1 == 5'h0; // @[RocketCore.scala 939:45]
  assign _T_765 = ibuf_io_inst_0_bits_inst_rs1; // @[RocketCore.scala 933:44]
  assign _T_768 = _T_760__T_767_data; // @[RocketCore.scala 939:25]
  assign _T_773 = ibuf_io_inst_0_bits_inst_rs2; // @[RocketCore.scala 933:44]
  assign _T_776 = _T_760__T_775_data; // @[RocketCore.scala 939:25]
  assign _T_847 = id_ctrl_csr == 3'h6; // @[package.scala 14:47]
  assign _T_848 = id_ctrl_csr == 3'h7; // @[package.scala 14:47]
  assign _T_849 = id_ctrl_csr == 3'h5; // @[package.scala 14:47]
  assign _T_850 = _T_847 | _T_848; // @[package.scala 14:62]
  assign id_csr_en = _T_850 | _T_849; // @[package.scala 14:62]
  assign id_system_insn = id_ctrl_csr == 3'h4; // @[RocketCore.scala 259:36]
  assign id_csr_ren = _T_850 & _T_763; // @[RocketCore.scala 260:54]
  assign _T_855 = id_ctrl_mem_cmd == 5'h14; // @[RocketCore.scala 262:50]
  assign id_sfence = id_ctrl_mem & _T_855; // @[RocketCore.scala 262:31]
  assign _T_856 = id_sfence | id_system_insn; // @[RocketCore.scala 263:32]
  assign _T_858 = id_csr_en & ~id_csr_ren; // @[RocketCore.scala 263:64]
  assign _T_859 = _T_858 & csr_io_decode_0_write_flush; // @[RocketCore.scala 263:79]
  assign id_csr_flush = _T_856 | _T_859; // @[RocketCore.scala 263:50]
  assign _T_864 = id_ctrl_div & ~csr_io_status_isa[12]; // @[RocketCore.scala 281:34]
  assign _T_865 = ~id_ctrl_legal | _T_864; // @[RocketCore.scala 280:40]
  assign _T_868 = id_ctrl_amo & ~csr_io_status_isa[0]; // @[RocketCore.scala 282:17]
  assign _T_869 = _T_865 | _T_868; // @[RocketCore.scala 281:65]
  assign _T_870 = csr_io_decode_0_fp_illegal | io_fpu_illegal_rm; // @[RocketCore.scala 283:48]
  assign _T_871 = id_ctrl_fp & _T_870; // @[RocketCore.scala 283:16]
  assign _T_872 = _T_869 | _T_871; // @[RocketCore.scala 282:48]
  assign _T_875 = id_ctrl_dp & ~csr_io_status_isa[3]; // @[RocketCore.scala 284:16]
  assign _T_876 = _T_872 | _T_875; // @[RocketCore.scala 283:70]
  assign _T_879 = ibuf_io_inst_0_bits_rvc & ~csr_io_status_isa[2]; // @[RocketCore.scala 285:30]
  assign _T_880 = _T_876 | _T_879; // @[RocketCore.scala 284:47]
  assign _T_886 = ~id_csr_ren & csr_io_decode_0_write_illegal; // @[RocketCore.scala 288:64]
  assign _T_887 = csr_io_decode_0_read_illegal | _T_886; // @[RocketCore.scala 288:49]
  assign _T_888 = id_csr_en & _T_887; // @[RocketCore.scala 288:15]
  assign _T_889 = _T_880 | _T_888; // @[RocketCore.scala 287:73]
  assign _T_892 = _T_856 & csr_io_decode_0_system_illegal; // @[RocketCore.scala 289:65]
  assign _T_893 = ~ibuf_io_inst_0_bits_rvc & _T_892; // @[RocketCore.scala 289:31]
  assign id_illegal_insn = _T_889 | _T_893; // @[RocketCore.scala 288:99]
  assign id_amo_aq = ibuf_io_inst_0_bits_inst_bits[26]; // @[RocketCore.scala 291:29]
  assign id_amo_rl = ibuf_io_inst_0_bits_inst_bits[25]; // @[RocketCore.scala 292:29]
  assign _T_894 = id_ctrl_amo & id_amo_aq; // @[RocketCore.scala 293:52]
  assign id_fence_next = id_ctrl_fence | _T_894; // @[RocketCore.scala 293:37]
  assign id_mem_busy = ~io_dmem_ordered | io_dmem_req_valid; // @[RocketCore.scala 294:38]
  assign _GEN_0 = id_mem_busy ? id_reg_fence : 1'h0; // @[RocketCore.scala 295:23]
  assign _T_904 = id_ctrl_amo & id_amo_rl; // @[RocketCore.scala 300:33]
  assign _T_905 = _T_904 | id_ctrl_fence_i; // @[RocketCore.scala 300:46]
  assign _T_907 = id_reg_fence & id_ctrl_mem; // @[RocketCore.scala 300:81]
  assign _T_908 = _T_905 | _T_907; // @[RocketCore.scala 300:65]
  assign id_do_fence = id_mem_busy & _T_908; // @[RocketCore.scala 300:17]
  assign _T_912 = csr_io_interrupt | bpu_io_debug_if; // @[RocketCore.scala 892:26]
  assign _T_913 = _T_912 | bpu_io_xcpt_if; // @[RocketCore.scala 892:26]
  assign _T_914 = _T_913 | ibuf_io_inst_0_bits_xcpt0_pf_inst; // @[RocketCore.scala 892:26]
  assign _T_915 = _T_914 | ibuf_io_inst_0_bits_xcpt0_ae_inst; // @[RocketCore.scala 892:26]
  assign _T_916 = _T_915 | ibuf_io_inst_0_bits_xcpt1_pf_inst; // @[RocketCore.scala 892:26]
  assign _T_917 = _T_916 | ibuf_io_inst_0_bits_xcpt1_ae_inst; // @[RocketCore.scala 892:26]
  assign id_xcpt = _T_917 | id_illegal_insn; // @[RocketCore.scala 892:26]
  assign _T_918 = ibuf_io_inst_0_bits_xcpt1_ae_inst ? 2'h1 : 2'h2; // @[Mux.scala 31:69]
  assign _T_919 = ibuf_io_inst_0_bits_xcpt1_pf_inst ? 4'hc : {{2'd0}, _T_918}; // @[Mux.scala 31:69]
  assign _T_920 = ibuf_io_inst_0_bits_xcpt0_ae_inst ? 4'h1 : _T_919; // @[Mux.scala 31:69]
  assign _T_921 = ibuf_io_inst_0_bits_xcpt0_pf_inst ? 4'hc : _T_920; // @[Mux.scala 31:69]
  assign _T_922 = bpu_io_xcpt_if ? 4'h3 : _T_921; // @[Mux.scala 31:69]
  assign _T_923 = bpu_io_debug_if ? 4'he : _T_922; // @[Mux.scala 31:69]
  assign ex_waddr = ex_reg_inst[11:7]; // @[RocketCore.scala 335:29]
  assign mem_waddr = mem_reg_inst[11:7]; // @[RocketCore.scala 336:31]
  assign wb_waddr = wb_reg_inst[11:7]; // @[RocketCore.scala 337:29]
  assign _T_934 = ex_reg_valid & ex_ctrl_wxd; // @[RocketCore.scala 340:19]
  assign _T_935 = mem_reg_valid & mem_ctrl_wxd; // @[RocketCore.scala 341:20]
  assign _T_937 = _T_935 & ~mem_ctrl_mem; // @[RocketCore.scala 341:36]
  assign _T_939 = 5'h0 == ibuf_io_inst_0_bits_inst_rs1; // @[RocketCore.scala 343:82]
  assign _T_941 = ex_waddr == ibuf_io_inst_0_bits_inst_rs1; // @[RocketCore.scala 343:82]
  assign _T_942 = _T_934 & _T_941; // @[RocketCore.scala 343:74]
  assign _T_943 = mem_waddr == ibuf_io_inst_0_bits_inst_rs1; // @[RocketCore.scala 343:82]
  assign _T_944 = _T_937 & _T_943; // @[RocketCore.scala 343:74]
  assign _T_946 = _T_935 & _T_943; // @[RocketCore.scala 343:74]
  assign _T_947 = 5'h0 == ibuf_io_inst_0_bits_inst_rs2; // @[RocketCore.scala 343:82]
  assign _T_949 = ex_waddr == ibuf_io_inst_0_bits_inst_rs2; // @[RocketCore.scala 343:82]
  assign _T_950 = _T_934 & _T_949; // @[RocketCore.scala 343:74]
  assign _T_951 = mem_waddr == ibuf_io_inst_0_bits_inst_rs2; // @[RocketCore.scala 343:82]
  assign _T_952 = _T_937 & _T_951; // @[RocketCore.scala 343:74]
  assign _T_954 = _T_935 & _T_951; // @[RocketCore.scala 343:74]
  assign _T_976 = ex_reg_rs_lsb_0 == 2'h1; // @[package.scala 31:81]
  assign _T_977 = _T_976 ? mem_reg_wdata : 64'h0; // @[package.scala 31:71]
  assign _T_978 = ex_reg_rs_lsb_0 == 2'h2; // @[package.scala 31:81]
  assign _T_979 = _T_978 ? wb_reg_wdata : _T_977; // @[package.scala 31:71]
  assign _T_980 = ex_reg_rs_lsb_0 == 2'h3; // @[package.scala 31:81]
  assign _T_981 = _T_980 ? io_dmem_resp_bits_data_word_bypass : _T_979; // @[package.scala 31:71]
  assign _T_982 = {ex_reg_rs_msb_0,ex_reg_rs_lsb_0}; // @[Cat.scala 30:58]
  assign _T_984 = ex_reg_rs_lsb_1 == 2'h1; // @[package.scala 31:81]
  assign _T_985 = _T_984 ? mem_reg_wdata : 64'h0; // @[package.scala 31:71]
  assign _T_986 = ex_reg_rs_lsb_1 == 2'h2; // @[package.scala 31:81]
  assign _T_987 = _T_986 ? wb_reg_wdata : _T_985; // @[package.scala 31:71]
  assign _T_988 = ex_reg_rs_lsb_1 == 2'h3; // @[package.scala 31:81]
  assign _T_989 = _T_988 ? io_dmem_resp_bits_data_word_bypass : _T_987; // @[package.scala 31:71]
  assign _T_990 = {ex_reg_rs_msb_1,ex_reg_rs_lsb_1}; // @[Cat.scala 30:58]
  assign _T_991 = ex_reg_rs_bypass_1 ? _T_989 : _T_990; // @[RocketCore.scala 351:14]
  assign _T_992 = ex_ctrl_sel_imm == 3'h5; // @[RocketCore.scala 954:24]
  assign _T_994 = ex_reg_inst[31]; // @[RocketCore.scala 954:53]
  assign _T_995 = _T_992 ? $signed(1'sh0) : $signed(_T_994); // @[RocketCore.scala 954:19]
  assign _T_996 = ex_ctrl_sel_imm == 3'h2; // @[RocketCore.scala 955:26]
  assign _T_998 = ex_reg_inst[30:20]; // @[RocketCore.scala 955:49]
  assign _T_1000 = ex_ctrl_sel_imm != 3'h2; // @[RocketCore.scala 956:26]
  assign _T_1001 = ex_ctrl_sel_imm != 3'h3; // @[RocketCore.scala 956:43]
  assign _T_1002 = _T_1000 & _T_1001; // @[RocketCore.scala 956:36]
  assign _T_1004 = ex_reg_inst[19:12]; // @[RocketCore.scala 956:73]
  assign _T_1008 = _T_996 | _T_992; // @[RocketCore.scala 957:33]
  assign _T_1009 = ex_ctrl_sel_imm == 3'h3; // @[RocketCore.scala 958:23]
  assign _T_1011 = ex_reg_inst[20]; // @[RocketCore.scala 958:44]
  assign _T_1012 = ex_ctrl_sel_imm == 3'h1; // @[RocketCore.scala 959:23]
  assign _T_1014 = ex_reg_inst[7]; // @[RocketCore.scala 959:43]
  assign _T_1015 = _T_1012 ? $signed(_T_1014) : $signed(_T_995); // @[RocketCore.scala 959:18]
  assign _T_1016 = _T_1009 ? $signed(_T_1011) : $signed(_T_1015); // @[RocketCore.scala 958:18]
  assign _T_1022 = _T_1008 ? 6'h0 : ex_reg_inst[30:25]; // @[RocketCore.scala 960:20]
  assign _T_1024 = ex_ctrl_sel_imm == 3'h0; // @[RocketCore.scala 962:24]
  assign _T_1026 = _T_1024 | _T_1012; // @[RocketCore.scala 962:34]
  assign _T_1031 = _T_992 ? ex_reg_inst[19:16] : ex_reg_inst[24:21]; // @[RocketCore.scala 963:19]
  assign _T_1032 = _T_1026 ? ex_reg_inst[11:8] : _T_1031; // @[RocketCore.scala 962:19]
  assign _T_1033 = _T_996 ? 4'h0 : _T_1032; // @[RocketCore.scala 961:19]
  assign _T_1036 = ex_ctrl_sel_imm == 3'h4; // @[RocketCore.scala 965:22]
  assign _T_1040 = _T_992 & ex_reg_inst[15]; // @[RocketCore.scala 966:17]
  assign _T_1041 = _T_1036 ? ex_reg_inst[20] : _T_1040; // @[RocketCore.scala 965:17]
  assign _T_1042 = _T_1024 ? ex_reg_inst[7] : _T_1041; // @[RocketCore.scala 964:17]
  assign _T_1045 = _T_1008 ? $signed(1'sh0) : $signed(_T_1016); // @[Cat.scala 30:58]
  assign _T_1046 = _T_1002 ? $signed({8{_T_995}}) : $signed(_T_1004); // @[Cat.scala 30:58]
  assign _T_1048 = _T_996 ? $signed(_T_998) : $signed({11{_T_995}}); // @[Cat.scala 30:58]
  assign _T_1049 = _T_992 ? $signed(1'sh0) : $signed(_T_994); // @[Cat.scala 30:58]
  assign ex_imm = {_T_1049,_T_1048,_T_1046,_T_1045,_T_1022,_T_1033,_T_1042}; // @[RocketCore.scala 968:53]
  assign _T_1053 = ex_reg_rs_bypass_0 ? _T_981 : _T_982; // @[RocketCore.scala 354:24]
  assign _T_1055 = 2'h2 == ex_ctrl_sel_alu1; // @[Mux.scala 46:19]
  assign _T_1056 = _T_1055 ? $signed(ex_reg_pc) : $signed(40'sh0); // @[Mux.scala 46:16]
  assign _T_1057 = 2'h1 == ex_ctrl_sel_alu1; // @[Mux.scala 46:19]
  assign _T_1058 = ex_reg_rs_bypass_1 ? _T_989 : _T_990; // @[RocketCore.scala 357:24]
  assign _T_1059 = ex_reg_rvc ? $signed(4'sh2) : $signed(4'sh4); // @[RocketCore.scala 359:19]
  assign _T_1060 = 2'h1 == ex_ctrl_sel_alu2; // @[Mux.scala 46:19]
  assign _T_1061 = _T_1060 ? $signed(_T_1059) : $signed(4'sh0); // @[Mux.scala 46:16]
  assign _T_1062 = 2'h3 == ex_ctrl_sel_alu2; // @[Mux.scala 46:19]
  assign _T_1063 = _T_1062 ? $signed(ex_imm) : $signed({{28{_T_1061[3]}},_T_1061}); // @[Mux.scala 46:16]
  assign _T_1064 = 2'h2 == ex_ctrl_sel_alu2; // @[Mux.scala 46:19]
  assign _T_1739 = ~ibuf_io_inst_0_valid | ibuf_io_inst_0_bits_replay; // @[RocketCore.scala 724:40]
  assign _T_1740 = _T_1739 | take_pc_mem_wb; // @[RocketCore.scala 724:71]
  assign _T_1543 = ibuf_io_inst_0_bits_inst_rs1 != 5'h0; // @[RocketCore.scala 656:55]
  assign _T_1544 = id_ctrl_rxs1 & _T_1543; // @[RocketCore.scala 656:42]
  assign _T_1591 = ibuf_io_inst_0_bits_inst_rs1 == ex_waddr; // @[RocketCore.scala 676:70]
  assign _T_1592 = _T_1544 & _T_1591; // @[RocketCore.scala 901:27]
  assign _T_1545 = ibuf_io_inst_0_bits_inst_rs2 != 5'h0; // @[RocketCore.scala 657:55]
  assign _T_1546 = id_ctrl_rxs2 & _T_1545; // @[RocketCore.scala 657:42]
  assign _T_1593 = ibuf_io_inst_0_bits_inst_rs2 == ex_waddr; // @[RocketCore.scala 676:70]
  assign _T_1594 = _T_1546 & _T_1593; // @[RocketCore.scala 901:27]
  assign _T_1597 = _T_1592 | _T_1594; // @[RocketCore.scala 901:50]
  assign _T_1547 = ibuf_io_inst_0_bits_inst_rd != 5'h0; // @[RocketCore.scala 658:55]
  assign _T_1548 = id_ctrl_wxd & _T_1547; // @[RocketCore.scala 658:42]
  assign _T_1595 = ibuf_io_inst_0_bits_inst_rd == ex_waddr; // @[RocketCore.scala 676:70]
  assign _T_1596 = _T_1548 & _T_1595; // @[RocketCore.scala 901:27]
  assign _T_1598 = _T_1597 | _T_1596; // @[RocketCore.scala 901:50]
  assign data_hazard_ex = ex_ctrl_wxd & _T_1598; // @[RocketCore.scala 676:36]
  assign _T_1585 = ex_ctrl_csr != 3'h0; // @[RocketCore.scala 675:38]
  assign _T_1586 = _T_1585 | ex_ctrl_jalr; // @[RocketCore.scala 675:48]
  assign _T_1587 = _T_1586 | ex_ctrl_mem; // @[RocketCore.scala 675:64]
  assign _T_1589 = _T_1587 | ex_ctrl_div; // @[RocketCore.scala 675:94]
  assign ex_cannot_bypass = _T_1589 | ex_ctrl_fp; // @[RocketCore.scala 675:109]
  assign _T_1610 = data_hazard_ex & ex_cannot_bypass; // @[RocketCore.scala 678:54]
  assign _T_1600 = io_fpu_dec_ren1 & _T_1591; // @[RocketCore.scala 901:27]
  assign _T_1602 = io_fpu_dec_ren2 & _T_1593; // @[RocketCore.scala 901:27]
  assign _T_1607 = _T_1600 | _T_1602; // @[RocketCore.scala 901:50]
  assign _T_1603 = ibuf_io_inst_0_bits_inst_rs3 == ex_waddr; // @[RocketCore.scala 677:76]
  assign _T_1604 = io_fpu_dec_ren3 & _T_1603; // @[RocketCore.scala 901:27]
  assign _T_1608 = _T_1607 | _T_1604; // @[RocketCore.scala 901:50]
  assign _T_1606 = io_fpu_dec_wen & _T_1595; // @[RocketCore.scala 901:27]
  assign _T_1609 = _T_1608 | _T_1606; // @[RocketCore.scala 901:50]
  assign fp_data_hazard_ex = ex_ctrl_wfd & _T_1609; // @[RocketCore.scala 677:39]
  assign _T_1611 = _T_1610 | fp_data_hazard_ex; // @[RocketCore.scala 678:74]
  assign id_ex_hazard = ex_reg_valid & _T_1611; // @[RocketCore.scala 678:35]
  assign _T_1618 = ibuf_io_inst_0_bits_inst_rs1 == mem_waddr; // @[RocketCore.scala 685:72]
  assign _T_1619 = _T_1544 & _T_1618; // @[RocketCore.scala 901:27]
  assign _T_1620 = ibuf_io_inst_0_bits_inst_rs2 == mem_waddr; // @[RocketCore.scala 685:72]
  assign _T_1621 = _T_1546 & _T_1620; // @[RocketCore.scala 901:27]
  assign _T_1624 = _T_1619 | _T_1621; // @[RocketCore.scala 901:50]
  assign _T_1622 = ibuf_io_inst_0_bits_inst_rd == mem_waddr; // @[RocketCore.scala 685:72]
  assign _T_1623 = _T_1548 & _T_1622; // @[RocketCore.scala 901:27]
  assign _T_1625 = _T_1624 | _T_1623; // @[RocketCore.scala 901:50]
  assign data_hazard_mem = mem_ctrl_wxd & _T_1625; // @[RocketCore.scala 685:38]
  assign _T_1612 = mem_ctrl_csr != 3'h0; // @[RocketCore.scala 684:40]
  assign _T_1613 = mem_ctrl_mem & mem_reg_slow_bypass; // @[RocketCore.scala 684:66]
  assign _T_1614 = _T_1612 | _T_1613; // @[RocketCore.scala 684:50]
  assign _T_1616 = _T_1614 | mem_ctrl_div; // @[RocketCore.scala 684:100]
  assign mem_cannot_bypass = _T_1616 | mem_ctrl_fp; // @[RocketCore.scala 684:116]
  assign _T_1637 = data_hazard_mem & mem_cannot_bypass; // @[RocketCore.scala 687:57]
  assign _T_1627 = io_fpu_dec_ren1 & _T_1618; // @[RocketCore.scala 901:27]
  assign _T_1629 = io_fpu_dec_ren2 & _T_1620; // @[RocketCore.scala 901:27]
  assign _T_1634 = _T_1627 | _T_1629; // @[RocketCore.scala 901:50]
  assign _T_1630 = ibuf_io_inst_0_bits_inst_rs3 == mem_waddr; // @[RocketCore.scala 686:78]
  assign _T_1631 = io_fpu_dec_ren3 & _T_1630; // @[RocketCore.scala 901:27]
  assign _T_1635 = _T_1634 | _T_1631; // @[RocketCore.scala 901:50]
  assign _T_1633 = io_fpu_dec_wen & _T_1622; // @[RocketCore.scala 901:27]
  assign _T_1636 = _T_1635 | _T_1633; // @[RocketCore.scala 901:50]
  assign fp_data_hazard_mem = mem_ctrl_wfd & _T_1636; // @[RocketCore.scala 686:41]
  assign _T_1638 = _T_1637 | fp_data_hazard_mem; // @[RocketCore.scala 687:78]
  assign id_mem_hazard = mem_reg_valid & _T_1638; // @[RocketCore.scala 687:37]
  assign _T_1711 = id_ex_hazard | id_mem_hazard; // @[RocketCore.scala 714:18]
  assign _T_1641 = ibuf_io_inst_0_bits_inst_rs1 == wb_waddr; // @[RocketCore.scala 691:70]
  assign _T_1642 = _T_1544 & _T_1641; // @[RocketCore.scala 901:27]
  assign _T_1643 = ibuf_io_inst_0_bits_inst_rs2 == wb_waddr; // @[RocketCore.scala 691:70]
  assign _T_1644 = _T_1546 & _T_1643; // @[RocketCore.scala 901:27]
  assign _T_1647 = _T_1642 | _T_1644; // @[RocketCore.scala 901:50]
  assign _T_1645 = ibuf_io_inst_0_bits_inst_rd == wb_waddr; // @[RocketCore.scala 691:70]
  assign _T_1646 = _T_1548 & _T_1645; // @[RocketCore.scala 901:27]
  assign _T_1648 = _T_1647 | _T_1646; // @[RocketCore.scala 901:50]
  assign data_hazard_wb = wb_ctrl_wxd & _T_1648; // @[RocketCore.scala 691:36]
  assign wb_dcache_miss = wb_ctrl_mem & ~io_dmem_resp_valid; // @[RocketCore.scala 448:36]
  assign wb_set_sboard = wb_ctrl_div | wb_dcache_miss; // @[RocketCore.scala 584:35]
  assign _T_1660 = data_hazard_wb & wb_set_sboard; // @[RocketCore.scala 693:54]
  assign _T_1650 = io_fpu_dec_ren1 & _T_1641; // @[RocketCore.scala 901:27]
  assign _T_1652 = io_fpu_dec_ren2 & _T_1643; // @[RocketCore.scala 901:27]
  assign _T_1657 = _T_1650 | _T_1652; // @[RocketCore.scala 901:50]
  assign _T_1653 = ibuf_io_inst_0_bits_inst_rs3 == wb_waddr; // @[RocketCore.scala 692:76]
  assign _T_1654 = io_fpu_dec_ren3 & _T_1653; // @[RocketCore.scala 901:27]
  assign _T_1658 = _T_1657 | _T_1654; // @[RocketCore.scala 901:50]
  assign _T_1656 = io_fpu_dec_wen & _T_1645; // @[RocketCore.scala 901:27]
  assign _T_1659 = _T_1658 | _T_1656; // @[RocketCore.scala 901:50]
  assign fp_data_hazard_wb = wb_ctrl_wfd & _T_1659; // @[RocketCore.scala 692:39]
  assign _T_1661 = _T_1660 | fp_data_hazard_wb; // @[RocketCore.scala 693:71]
  assign id_wb_hazard = wb_reg_valid & _T_1661; // @[RocketCore.scala 693:35]
  assign _T_1712 = _T_1711 | id_wb_hazard; // @[RocketCore.scala 714:35]
  assign _T_1552 = {_T_1550[31:1], 1'h0}; // @[RocketCore.scala 919:40]
  assign _T_1558 = _T_1552 >> ibuf_io_inst_0_bits_inst_rs1; // @[RocketCore.scala 915:35]
  assign dmem_resp_valid = io_dmem_resp_valid & io_dmem_resp_bits_has_data; // @[RocketCore.scala 594:44]
  assign dmem_resp_replay = dmem_resp_valid & io_dmem_resp_bits_replay; // @[RocketCore.scala 595:42]
  assign dmem_resp_xpu = ~io_dmem_resp_bits_tag[0]; // @[RocketCore.scala 591:23]
  assign _T_1486 = dmem_resp_replay & dmem_resp_xpu; // @[RocketCore.scala 610:26]
  assign _T_1484 = div_io_resp_ready & div_io_resp_valid; // @[Decoupled.scala 37:37]
  assign ll_wen = _T_1486 | _T_1484; // @[RocketCore.scala 610:44]
  assign dmem_resp_waddr = io_dmem_resp_bits_tag[5:1]; // @[RocketCore.scala 593:46]
  assign ll_waddr = _T_1486 ? dmem_resp_waddr : div_io_resp_bits_tag; // @[RocketCore.scala 610:44]
  assign _T_1560 = ll_waddr == ibuf_io_inst_0_bits_inst_rs1; // @[RocketCore.scala 668:70]
  assign _T_1561 = ll_wen & _T_1560; // @[RocketCore.scala 668:58]
  assign _T_1563 = _T_1558[0] & ~_T_1561; // @[RocketCore.scala 671:77]
  assign _T_1564 = _T_1544 & _T_1563; // @[RocketCore.scala 901:27]
  assign _T_1565 = _T_1552 >> ibuf_io_inst_0_bits_inst_rs2; // @[RocketCore.scala 915:35]
  assign _T_1567 = ll_waddr == ibuf_io_inst_0_bits_inst_rs2; // @[RocketCore.scala 668:70]
  assign _T_1568 = ll_wen & _T_1567; // @[RocketCore.scala 668:58]
  assign _T_1570 = _T_1565[0] & ~_T_1568; // @[RocketCore.scala 671:77]
  assign _T_1571 = _T_1546 & _T_1570; // @[RocketCore.scala 901:27]
  assign _T_1579 = _T_1564 | _T_1571; // @[RocketCore.scala 901:50]
  assign _T_1572 = _T_1552 >> ibuf_io_inst_0_bits_inst_rd; // @[RocketCore.scala 915:35]
  assign _T_1574 = ll_waddr == ibuf_io_inst_0_bits_inst_rd; // @[RocketCore.scala 668:70]
  assign _T_1575 = ll_wen & _T_1574; // @[RocketCore.scala 668:58]
  assign _T_1577 = _T_1572[0] & ~_T_1575; // @[RocketCore.scala 671:77]
  assign _T_1578 = _T_1548 & _T_1577; // @[RocketCore.scala 901:27]
  assign id_sboard_hazard = _T_1579 | _T_1578; // @[RocketCore.scala 901:50]
  assign _T_1713 = _T_1712 | id_sboard_hazard; // @[RocketCore.scala 714:51]
  assign _T_1714 = ex_reg_valid | mem_reg_valid; // @[RocketCore.scala 715:40]
  assign _T_1715 = _T_1714 | wb_reg_valid; // @[RocketCore.scala 715:57]
  assign _T_1716 = csr_io_singleStep & _T_1715; // @[RocketCore.scala 715:23]
  assign _T_1717 = _T_1713 | _T_1716; // @[RocketCore.scala 714:71]
  assign _T_1718 = id_csr_en & csr_io_decode_0_fp_csr; // @[RocketCore.scala 716:15]
  assign _T_1720 = _T_1718 & ~io_fpu_fcsr_rdy; // @[RocketCore.scala 716:42]
  assign _T_1721 = _T_1717 | _T_1720; // @[RocketCore.scala 715:74]
  assign _T_1682 = _T_1663 >> ibuf_io_inst_0_bits_inst_rs1; // @[RocketCore.scala 915:35]
  assign _T_1684 = io_fpu_dec_ren1 & _T_1682[0]; // @[RocketCore.scala 901:27]
  assign _T_1685 = _T_1663 >> ibuf_io_inst_0_bits_inst_rs2; // @[RocketCore.scala 915:35]
  assign _T_1687 = io_fpu_dec_ren2 & _T_1685[0]; // @[RocketCore.scala 901:27]
  assign _T_1694 = _T_1684 | _T_1687; // @[RocketCore.scala 901:50]
  assign _T_1688 = _T_1663 >> ibuf_io_inst_0_bits_inst_rs3; // @[RocketCore.scala 915:35]
  assign _T_1690 = io_fpu_dec_ren3 & _T_1688[0]; // @[RocketCore.scala 901:27]
  assign _T_1695 = _T_1694 | _T_1690; // @[RocketCore.scala 901:50]
  assign _T_1691 = _T_1663 >> ibuf_io_inst_0_bits_inst_rd; // @[RocketCore.scala 915:35]
  assign _T_1693 = io_fpu_dec_wen & _T_1691[0]; // @[RocketCore.scala 901:27]
  assign id_stall_fpu = _T_1695 | _T_1693; // @[RocketCore.scala 901:50]
  assign _T_1722 = id_ctrl_fp & id_stall_fpu; // @[RocketCore.scala 717:16]
  assign _T_1723 = _T_1721 | _T_1722; // @[RocketCore.scala 716:62]
  assign dcache_blocked = blocked & ~io_dmem_perf_grant; // @[RocketCore.scala 708:13]
  assign _T_1724 = id_ctrl_mem & dcache_blocked; // @[RocketCore.scala 718:17]
  assign _T_1725 = _T_1723 | _T_1724; // @[RocketCore.scala 717:32]
  assign wb_wxd = wb_reg_valid & wb_ctrl_wxd; // @[RocketCore.scala 583:29]
  assign _T_1729 = div_io_resp_valid & ~wb_wxd; // @[RocketCore.scala 720:62]
  assign _T_1730 = div_io_req_ready | _T_1729; // @[RocketCore.scala 720:40]
  assign _T_1732 = ~_T_1730 | div_io_req_valid; // @[RocketCore.scala 720:75]
  assign _T_1733 = id_ctrl_div & _T_1732; // @[RocketCore.scala 720:17]
  assign _T_1734 = _T_1725 | _T_1733; // @[RocketCore.scala 719:34]
  assign _T_1737 = _T_1734 | id_do_fence; // @[RocketCore.scala 721:15]
  assign ctrl_stalld = _T_1737 | csr_io_csr_stall; // @[RocketCore.scala 722:17]
  assign _T_1741 = _T_1740 | ctrl_stalld; // @[RocketCore.scala 724:89]
  assign ctrl_killd = _T_1741 | csr_io_interrupt; // @[RocketCore.scala 724:104]
  assign _T_1070 = ~take_pc_mem_wb & ibuf_io_inst_0_valid; // @[RocketCore.scala 391:29]
  assign _GEN_1 = id_fence_next | _GEN_0; // @[RocketCore.scala 399:26]
  assign _T_1078 = {ibuf_io_inst_0_bits_xcpt1_pf_inst,ibuf_io_inst_0_bits_xcpt1_ae_inst}; // @[RocketCore.scala 405:22]
  assign _T_1079 = _T_1078 != 2'h0; // @[RocketCore.scala 405:29]
  assign _GEN_4 = _T_1079 | ibuf_io_inst_0_bits_rvc; // @[RocketCore.scala 405:34]
  assign _T_1080 = {ibuf_io_inst_0_bits_xcpt0_pf_inst,ibuf_io_inst_0_bits_xcpt0_ae_inst}; // @[RocketCore.scala 410:40]
  assign _T_1081 = _T_1080 != 2'h0; // @[RocketCore.scala 410:47]
  assign _T_1082 = bpu_io_xcpt_if | _T_1081; // @[RocketCore.scala 410:28]
  assign _GEN_8 = id_xcpt | id_ctrl_alu_dw; // @[RocketCore.scala 400:20]
  assign _T_1083 = id_ctrl_fence_i | id_csr_flush; // @[RocketCore.scala 415:42]
  assign _T_1086 = {_T_1545,_T_1543}; // @[Cat.scala 30:58]
  assign _T_1087 = _T_939 | _T_942; // @[RocketCore.scala 422:48]
  assign _T_1088 = _T_1087 | _T_944; // @[RocketCore.scala 422:48]
  assign do_bypass = _T_1088 | _T_946; // @[RocketCore.scala 422:48]
  assign _T_1092 = id_ctrl_rxs1 & ~do_bypass; // @[RocketCore.scala 426:23]
  assign _T_1488 = wb_reg_valid & ~replay_wb_common; // @[RocketCore.scala 618:31]
  assign wb_valid = _T_1488 & ~wb_xcpt; // @[RocketCore.scala 618:45]
  assign wb_wen = wb_valid & wb_ctrl_wxd; // @[RocketCore.scala 619:25]
  assign rf_wen = wb_wen | ll_wen; // @[RocketCore.scala 620:23]
  assign rf_waddr = ll_wen ? ll_waddr : wb_waddr; // @[RocketCore.scala 621:21]
  assign _T_1496 = rf_waddr != 5'h0; // @[RocketCore.scala 944:16]
  assign _T_1500 = rf_waddr == ibuf_io_inst_0_bits_inst_rs1; // @[RocketCore.scala 947:20]
  assign _T_1490 = dmem_resp_valid & dmem_resp_xpu; // @[RocketCore.scala 622:38]
  assign ll_wdata = div_io_resp_bits_data;
  assign _T_1492 = wb_ctrl_csr != 3'h0; // @[RocketCore.scala 624:34]
  assign _T_1494 = _T_1492 ? csr_io_rw_rdata : wb_reg_wdata; // @[RocketCore.scala 624:21]
  assign _T_1495 = ll_wen ? ll_wdata : _T_1494; // @[RocketCore.scala 623:21]
  assign rf_wdata = _T_1490 ? io_dmem_resp_bits_data : _T_1495; // @[RocketCore.scala 622:21]
  assign _GEN_214 = _T_1500 ? rf_wdata : _T_768; // @[RocketCore.scala 947:31]
  assign _GEN_221 = _T_1496 ? _GEN_214 : _T_768; // @[RocketCore.scala 944:29]
  assign _GEN_228 = rf_wen ? _GEN_221 : _T_768; // @[RocketCore.scala 627:17]
  assign _T_1095 = _T_947 | _T_950; // @[RocketCore.scala 422:48]
  assign _T_1096 = _T_1095 | _T_952; // @[RocketCore.scala 422:48]
  assign do_bypass_1 = _T_1096 | _T_954; // @[RocketCore.scala 422:48]
  assign _T_1100 = id_ctrl_rxs2 & ~do_bypass_1; // @[RocketCore.scala 426:23]
  assign _T_1501 = rf_waddr == ibuf_io_inst_0_bits_inst_rs2; // @[RocketCore.scala 947:20]
  assign _GEN_215 = _T_1501 ? rf_wdata : _T_776; // @[RocketCore.scala 947:31]
  assign _GEN_222 = _T_1496 ? _GEN_215 : _T_776; // @[RocketCore.scala 944:29]
  assign _GEN_229 = rf_wen ? _GEN_222 : _T_776; // @[RocketCore.scala 627:17]
  assign inst = ibuf_io_inst_0_bits_rvc ? {{16'd0}, ibuf_io_inst_0_bits_raw[15:0]} : ibuf_io_inst_0_bits_raw; // @[RocketCore.scala 432:21]
  assign _T_1639 = mem_reg_valid & data_hazard_mem; // @[RocketCore.scala 688:32]
  assign id_load_use = _T_1639 & mem_ctrl_mem; // @[RocketCore.scala 688:51]
  assign _T_1107 = ~ctrl_killd | csr_io_interrupt; // @[RocketCore.scala 438:21]
  assign _T_1108 = _T_1107 | ibuf_io_inst_0_bits_replay; // @[RocketCore.scala 438:41]
  assign _T_1112 = ex_ctrl_mem & ~io_dmem_req_ready; // @[RocketCore.scala 449:42]
  assign _T_1114 = ex_ctrl_div & ~div_io_req_ready; // @[RocketCore.scala 450:42]
  assign replay_ex_structural = _T_1112 | _T_1114; // @[RocketCore.scala 449:64]
  assign replay_ex_load_use = wb_dcache_miss & ex_reg_load_use; // @[RocketCore.scala 451:43]
  assign _T_1115 = replay_ex_structural | replay_ex_load_use; // @[RocketCore.scala 452:75]
  assign _T_1116 = ex_reg_valid & _T_1115; // @[RocketCore.scala 452:50]
  assign replay_ex = ex_reg_replay | _T_1116; // @[RocketCore.scala 452:33]
  assign _T_1117 = take_pc_mem_wb | replay_ex; // @[RocketCore.scala 453:35]
  assign ctrl_killx = _T_1117 | ~ex_reg_valid; // @[RocketCore.scala 453:48]
  assign _T_1119 = ex_ctrl_mem_cmd == 5'h7; // @[RocketCore.scala 455:40]
  assign _T_1130 = 3'h0 == ex_ctrl_mem_type; // @[RocketCore.scala 455:91]
  assign _T_1131 = 3'h4 == ex_ctrl_mem_type; // @[RocketCore.scala 455:91]
  assign _T_1132 = 3'h1 == ex_ctrl_mem_type; // @[RocketCore.scala 455:91]
  assign _T_1133 = 3'h5 == ex_ctrl_mem_type; // @[RocketCore.scala 455:91]
  assign _T_1135 = _T_1130 | _T_1131; // @[RocketCore.scala 455:91]
  assign _T_1136 = _T_1135 | _T_1132; // @[RocketCore.scala 455:91]
  assign _T_1137 = _T_1136 | _T_1133; // @[RocketCore.scala 455:91]
  assign ex_slow_bypass = _T_1119 | _T_1137; // @[RocketCore.scala 455:50]
  assign _T_1139 = ex_ctrl_mem_cmd == 5'h14; // @[RocketCore.scala 456:67]
  assign ex_sfence = ex_ctrl_mem & _T_1139; // @[RocketCore.scala 456:48]
  assign ex_xcpt = ex_reg_xcpt_interrupt | ex_reg_xcpt; // @[RocketCore.scala 459:28]
  assign _T_1150 = mem_reg_valid | mem_reg_replay; // @[RocketCore.scala 465:36]
  assign mem_pc_valid = _T_1150 | mem_reg_xcpt_interrupt; // @[RocketCore.scala 465:54]
  assign _T_1303 = ~csr_io_status_isa[2] & mem_npc[1]; // @[RocketCore.scala 474:56]
  assign mem_npc_misaligned = _T_1303 & ~mem_reg_sfence; // @[RocketCore.scala 474:70]
  assign _T_1306 = mem_ctrl_jalr ^ mem_npc_misaligned; // @[RocketCore.scala 475:59]
  assign _T_1307 = ~mem_reg_xcpt & _T_1306; // @[RocketCore.scala 475:41]
  assign mem_int_wdata = _T_1307 ? $signed({{24{mem_br_target[39]}},mem_br_target}) : $signed(mem_reg_wdata); // @[RocketCore.scala 475:119]
  assign _T_1310 = mem_ctrl_branch | mem_ctrl_jalr; // @[RocketCore.scala 476:33]
  assign mem_cfi = _T_1310 | mem_ctrl_jal; // @[RocketCore.scala 476:50]
  assign _T_1312 = _T_1152 | mem_ctrl_jalr; // @[RocketCore.scala 477:57]
  assign mem_cfi_taken = _T_1312 | mem_ctrl_jal; // @[RocketCore.scala 477:74]
  assign _T_1324 = mem_reg_valid & mem_reg_flush_pipe; // @[RocketCore.scala 489:23]
  assign _T_1325 = ex_ctrl_mem_cmd == 5'h0; // @[Consts.scala 93:31]
  assign _T_1326 = ex_ctrl_mem_cmd == 5'h6; // @[Consts.scala 93:48]
  assign _T_1327 = _T_1325 | _T_1326; // @[Consts.scala 93:41]
  assign _T_1329 = _T_1327 | _T_1119; // @[Consts.scala 93:58]
  assign _T_1330 = ex_ctrl_mem_cmd == 5'h4; // @[package.scala 14:47]
  assign _T_1331 = ex_ctrl_mem_cmd == 5'h9; // @[package.scala 14:47]
  assign _T_1332 = ex_ctrl_mem_cmd == 5'ha; // @[package.scala 14:47]
  assign _T_1333 = ex_ctrl_mem_cmd == 5'hb; // @[package.scala 14:47]
  assign _T_1334 = _T_1330 | _T_1331; // @[package.scala 14:62]
  assign _T_1335 = _T_1334 | _T_1332; // @[package.scala 14:62]
  assign _T_1336 = _T_1335 | _T_1333; // @[package.scala 14:62]
  assign _T_1337 = ex_ctrl_mem_cmd == 5'h8; // @[package.scala 14:47]
  assign _T_1338 = ex_ctrl_mem_cmd == 5'hc; // @[package.scala 14:47]
  assign _T_1339 = ex_ctrl_mem_cmd == 5'hd; // @[package.scala 14:47]
  assign _T_1340 = ex_ctrl_mem_cmd == 5'he; // @[package.scala 14:47]
  assign _T_1341 = ex_ctrl_mem_cmd == 5'hf; // @[package.scala 14:47]
  assign _T_1342 = _T_1337 | _T_1338; // @[package.scala 14:62]
  assign _T_1343 = _T_1342 | _T_1339; // @[package.scala 14:62]
  assign _T_1344 = _T_1343 | _T_1340; // @[package.scala 14:62]
  assign _T_1345 = _T_1344 | _T_1341; // @[package.scala 14:62]
  assign _T_1346 = _T_1336 | _T_1345; // @[Consts.scala 91:44]
  assign _T_1347 = _T_1329 | _T_1346; // @[Consts.scala 93:75]
  assign _T_1348 = ex_ctrl_mem & _T_1347; // @[RocketCore.scala 494:33]
  assign _T_1349 = ex_ctrl_mem_cmd == 5'h1; // @[Consts.scala 94:32]
  assign _T_1350 = ex_ctrl_mem_cmd == 5'h11; // @[Consts.scala 94:49]
  assign _T_1351 = _T_1349 | _T_1350; // @[Consts.scala 94:42]
  assign _T_1353 = _T_1351 | _T_1119; // @[Consts.scala 94:59]
  assign _T_1371 = _T_1353 | _T_1346; // @[Consts.scala 94:76]
  assign _T_1372 = ex_ctrl_mem & _T_1371; // @[RocketCore.scala 495:34]
  assign _T_1374 = ex_ctrl_mem | ex_sfence; // @[RocketCore.scala 508:56]
  assign _T_1375 = ex_ctrl_rxs2 & _T_1374; // @[RocketCore.scala 508:24]
  assign _T_1377 = ex_ctrl_mem_type[1:0] == 2'h0; // @[AMOALU.scala 26:19]
  assign _T_1381 = {_T_991[7:0],_T_991[7:0],_T_991[7:0],_T_991[7:0],_T_991[7:0],_T_991[7:0],_T_991[7:0],_T_991[7:0]}; // @[Cat.scala 30:58]
  assign _T_1382 = ex_ctrl_mem_type[1:0] == 2'h1; // @[AMOALU.scala 26:19]
  assign _T_1385 = {_T_991[15:0],_T_991[15:0],_T_991[15:0],_T_991[15:0]}; // @[Cat.scala 30:58]
  assign _T_1386 = ex_ctrl_mem_type[1:0] == 2'h2; // @[AMOALU.scala 26:19]
  assign _T_1388 = {_T_991[31:0],_T_991[31:0]}; // @[Cat.scala 30:58]
  assign _T_1392 = ex_ctrl_jalr & csr_io_status_debug; // @[RocketCore.scala 512:24]
  assign _GEN_72 = _T_1392 | ex_ctrl_fence_i; // @[RocketCore.scala 512:48]
  assign _GEN_73 = _T_1392 | ex_reg_flush_pipe; // @[RocketCore.scala 512:48]
  assign _T_1393 = mem_reg_load & bpu_io_xcpt_ld; // @[RocketCore.scala 519:38]
  assign _T_1394 = mem_reg_store & bpu_io_xcpt_st; // @[RocketCore.scala 519:75]
  assign mem_breakpoint = _T_1393 | _T_1394; // @[RocketCore.scala 519:57]
  assign _T_1395 = mem_reg_load & bpu_io_debug_ld; // @[RocketCore.scala 520:44]
  assign _T_1396 = mem_reg_store & bpu_io_debug_st; // @[RocketCore.scala 520:82]
  assign mem_debug_breakpoint = _T_1395 | _T_1396; // @[RocketCore.scala 520:64]
  assign mem_ldst_xcpt = mem_debug_breakpoint | mem_breakpoint; // @[RocketCore.scala 892:26]
  assign mem_ldst_cause = mem_debug_breakpoint ? 4'he : 4'h3; // @[Mux.scala 31:69]
  assign _T_1397 = mem_reg_xcpt_interrupt | mem_reg_xcpt; // @[RocketCore.scala 526:29]
  assign _T_1398 = mem_reg_valid & mem_npc_misaligned; // @[RocketCore.scala 527:20]
  assign _T_1399 = mem_reg_valid & mem_ldst_xcpt; // @[RocketCore.scala 528:20]
  assign _T_1400 = _T_1397 | _T_1398; // @[RocketCore.scala 892:26]
  assign mem_xcpt = _T_1400 | _T_1399; // @[RocketCore.scala 892:26]
  assign _T_1401 = _T_1398 ? 4'h0 : mem_ldst_cause; // @[Mux.scala 31:69]
  assign dcache_kill_mem = _T_935 & io_dmem_replay_next; // @[RocketCore.scala 537:55]
  assign _T_1415 = mem_reg_valid & mem_ctrl_fp; // @[RocketCore.scala 538:36]
  assign fpu_kill_mem = _T_1415 & io_fpu_nack_mem; // @[RocketCore.scala 538:51]
  assign _T_1416 = dcache_kill_mem | mem_reg_replay; // @[RocketCore.scala 539:37]
  assign replay_mem = _T_1416 | fpu_kill_mem; // @[RocketCore.scala 539:55]
  assign _T_1417 = dcache_kill_mem | take_pc_wb; // @[RocketCore.scala 540:38]
  assign _T_1418 = _T_1417 | mem_reg_xcpt; // @[RocketCore.scala 540:52]
  assign killm_common = _T_1418 | ~mem_reg_valid; // @[RocketCore.scala 540:68]
  assign _T_1424 = killm_common | mem_xcpt; // @[RocketCore.scala 542:33]
  assign ctrl_killm = _T_1424 | fpu_kill_mem; // @[RocketCore.scala 542:45]
  assign _T_1433 = ~mem_reg_xcpt & mem_ctrl_fp; // @[RocketCore.scala 552:39]
  assign _T_1434 = _T_1433 & mem_ctrl_wxd; // @[RocketCore.scala 552:54]
  assign _T_1454 = _T_1446 ? 3'h7 : 3'h5; // @[Mux.scala 31:69]
  assign _T_1455 = _T_1444 ? 4'hd : {{1'd0}, _T_1454}; // @[Mux.scala 31:69]
  assign _T_1456 = _T_1442 ? 4'hf : _T_1455; // @[Mux.scala 31:69]
  assign _T_1457 = _T_1440 ? 4'h4 : _T_1456; // @[Mux.scala 31:69]
  assign _T_1458 = _T_1438 ? 4'h6 : _T_1457; // @[Mux.scala 31:69]
  assign wb_cause = wb_reg_xcpt ? wb_reg_cause : {{60'd0}, _T_1458}; // @[Mux.scala 31:69]
  assign _T_1459 = wb_cause == 64'h6; // @[RocketCore.scala 896:38]
  assign _T_1461 = wb_cause == 64'h4; // @[RocketCore.scala 896:38]
  assign _T_1463 = wb_cause == 64'hf; // @[RocketCore.scala 896:38]
  assign _T_1465 = wb_cause == 64'hd; // @[RocketCore.scala 896:38]
  assign _T_1467 = wb_cause == 64'h7; // @[RocketCore.scala 896:38]
  assign _T_1469 = wb_cause == 64'h5; // @[RocketCore.scala 896:38]
  assign _T_1510 = wb_cause == 64'h2; // @[package.scala 14:47]
  assign _T_1511 = wb_cause == 64'h3; // @[package.scala 14:47]
  assign _T_1516 = wb_cause == 64'h1; // @[package.scala 14:47]
  assign _T_1519 = wb_cause == 64'hc; // @[package.scala 14:47]
  assign _T_1520 = _T_1510 | _T_1511; // @[package.scala 14:62]
  assign _T_1521 = _T_1520 | _T_1461; // @[package.scala 14:62]
  assign _T_1522 = _T_1521 | _T_1459; // @[package.scala 14:62]
  assign _T_1523 = _T_1522 | _T_1469; // @[package.scala 14:62]
  assign _T_1524 = _T_1523 | _T_1467; // @[package.scala 14:62]
  assign _T_1525 = _T_1524 | _T_1516; // @[package.scala 14:62]
  assign _T_1526 = _T_1525 | _T_1465; // @[package.scala 14:62]
  assign _T_1527 = _T_1526 | _T_1463; // @[package.scala 14:62]
  assign _T_1528 = _T_1527 | _T_1519; // @[package.scala 14:62]
  assign tval_valid = wb_xcpt & _T_1528; // @[RocketCore.scala 642:28]
  assign a_1 = wb_reg_wdata[63:39]; // @[RocketCore.scala 906:23]
  assign _T_1530 = $signed(a_1) == 25'sh0; // @[RocketCore.scala 907:21]
  assign _T_1531 = $signed(a_1) == -25'sh1; // @[RocketCore.scala 907:34]
  assign _T_1532 = _T_1530 | _T_1531; // @[RocketCore.scala 907:29]
  assign msb_1 = _T_1532 ? wb_reg_wdata[39] : ~wb_reg_wdata[38]; // @[RocketCore.scala 907:18]
  assign _T_1537 = {msb_1,wb_reg_wdata[38:0]}; // @[Cat.scala 30:58]
  assign _T_1540 = wb_reg_valid ? 3'h0 : 3'h4; // @[CSR.scala 128:15]
  assign _T_1553 = 32'h1 << ll_waddr; // @[RocketCore.scala 922:62]
  assign _T_1554 = ll_wen ? _T_1553 : 32'h0; // @[RocketCore.scala 922:49]
  assign _T_1556 = _T_1552 & ~_T_1554; // @[RocketCore.scala 914:62]
  assign _T_1580 = wb_set_sboard & wb_wen; // @[RocketCore.scala 672:28]
  assign _T_1581 = 32'h1 << wb_waddr; // @[RocketCore.scala 922:62]
  assign _T_1582 = _T_1580 ? _T_1581 : 32'h0; // @[RocketCore.scala 922:49]
  assign _T_1583 = _T_1556 | _T_1582; // @[RocketCore.scala 913:60]
  assign _T_1584 = ll_wen | _T_1580; // @[RocketCore.scala 925:17]
  assign _T_1664 = wb_dcache_miss & wb_ctrl_wfd; // @[RocketCore.scala 697:35]
  assign _T_1665 = _T_1664 | io_fpu_sboard_set; // @[RocketCore.scala 697:50]
  assign _T_1666 = _T_1665 & wb_valid; // @[RocketCore.scala 697:72]
  assign _T_1668 = _T_1666 ? _T_1581 : 32'h0; // @[RocketCore.scala 922:49]
  assign _T_1669 = _T_1663 | _T_1668; // @[RocketCore.scala 913:60]
  assign _T_1671 = dmem_resp_replay & io_dmem_resp_bits_tag[0]; // @[RocketCore.scala 698:38]
  assign _T_1672 = 32'h1 << dmem_resp_waddr; // @[RocketCore.scala 922:62]
  assign _T_1673 = _T_1671 ? _T_1672 : 32'h0; // @[RocketCore.scala 922:49]
  assign _T_1675 = _T_1669 & ~_T_1673; // @[RocketCore.scala 914:62]
  assign _T_1676 = _T_1666 | _T_1671; // @[RocketCore.scala 925:17]
  assign _T_1677 = 32'h1 << io_fpu_sboard_clra; // @[RocketCore.scala 922:62]
  assign _T_1678 = io_fpu_sboard_clr ? _T_1677 : 32'h0; // @[RocketCore.scala 922:49]
  assign _T_1680 = _T_1675 & ~_T_1678; // @[RocketCore.scala 914:62]
  assign _T_1681 = _T_1676 | io_fpu_sboard_clr; // @[RocketCore.scala 925:17]
  assign _T_1698 = ~io_dmem_req_ready & io_dmem_clock_enabled; // @[RocketCore.scala 707:35]
  assign _T_1700 = _T_1698 & ~io_dmem_perf_grant; // @[RocketCore.scala 707:60]
  assign _T_1701 = blocked | io_dmem_req_valid; // @[RocketCore.scala 707:95]
  assign _T_1702 = _T_1701 | io_dmem_s2_nack; // @[RocketCore.scala 707:116]
  assign _T_1744 = wb_xcpt | csr_io_eret; // @[RocketCore.scala 729:17]
  assign _T_1745 = replay_wb_common ? wb_reg_pc : mem_npc; // @[RocketCore.scala 730:8]
  assign _T_1747 = wb_reg_valid & wb_ctrl_fence_i; // @[RocketCore.scala 732:40]
  assign _T_1750 = ex_pc_valid | mem_pc_valid; // @[RocketCore.scala 734:43]
  assign _T_1758 = mem_reg_valid & ~take_pc_wb; // @[RocketCore.scala 746:45]
  assign _T_1759 = _T_1758 & mem_wrong_npc; // @[RocketCore.scala 746:60]
  assign _T_1761 = ~mem_cfi | mem_cfi_taken; // @[RocketCore.scala 746:90]
  assign _T_1763 = mem_ctrl_jal | mem_ctrl_jalr; // @[RocketCore.scala 749:23]
  assign _T_1765 = _T_1763 & mem_waddr[0]; // @[RocketCore.scala 749:41]
  assign _T_1767 = mem_reg_inst[19:15] & 5'h1b; // @[RocketCore.scala 750:46]
  assign _T_1768 = 5'h1 == _T_1767; // @[RocketCore.scala 750:46]
  assign _T_1769 = mem_ctrl_jalr & _T_1768; // @[RocketCore.scala 750:23]
  assign _T_1772 = _T_1769 ? 2'h3 : {{1'd0}, _T_1763}; // @[RocketCore.scala 750:8]
  assign _T_1774 = mem_reg_rvc ? 2'h0 : 2'h2; // @[RocketCore.scala 754:74]
  assign _GEN_237 = {{38'd0}, _T_1774}; // @[RocketCore.scala 754:69]
  assign _T_1776 = mem_reg_pc + _GEN_237; // @[RocketCore.scala 754:69]
  assign _T_1778 = ~io_imem_btb_update_bits_br_pc | 39'h3; // @[RocketCore.scala 755:66]
  assign ex_dcache_tag = {ex_waddr,ex_ctrl_fp}; // @[Cat.scala 30:58]
  assign a_2 = _T_1053[63:39]; // @[RocketCore.scala 906:23]
  assign _T_1788 = $signed(a_2) == 25'sh0; // @[RocketCore.scala 907:21]
  assign _T_1789 = $signed(a_2) == -25'sh1; // @[RocketCore.scala 907:34]
  assign _T_1790 = _T_1788 | _T_1789; // @[RocketCore.scala 907:29]
  assign msb_2 = _T_1790 ? alu_io_adder_out[39] : ~alu_io_adder_out[38]; // @[RocketCore.scala 907:18]
  assign _T_1797 = killm_common | mem_ldst_xcpt; // @[RocketCore.scala 785:35]
  assign io_imem_might_request = imem_might_request_reg; // @[RocketCore.scala 733:25]
  assign io_imem_req_valid = take_pc_wb | take_pc_mem; // @[RocketCore.scala 726:21]
  assign io_imem_req_bits_pc = _T_1744 ? csr_io_evec : _T_1745; // @[RocketCore.scala 728:23]
  assign io_imem_req_bits_speculative = ~take_pc_wb; // @[RocketCore.scala 727:32]
  assign io_imem_sfence_valid = wb_reg_valid & wb_reg_sfence; // @[RocketCore.scala 737:24]
  assign io_imem_sfence_bits_rs1 = wb_ctrl_mem_type[0]; // @[RocketCore.scala 738:27]
  assign io_imem_sfence_bits_rs2 = wb_ctrl_mem_type[1]; // @[RocketCore.scala 739:27]
  assign io_imem_sfence_bits_addr = wb_reg_wdata[38:0]; // @[RocketCore.scala 740:28]
  assign io_imem_resp_ready = ibuf_io_imem_ready; // @[RocketCore.scala 240:16]
  assign io_imem_btb_update_valid = _T_1759 & _T_1761; // @[RocketCore.scala 746:28]
  assign io_imem_btb_update_bits_prediction_entry = mem_reg_btb_resp_entry; // @[RocketCore.scala 756:38]
  assign io_imem_btb_update_bits_pc = ~_T_1778; // @[RocketCore.scala 755:30]
  assign io_imem_btb_update_bits_isValid = _T_1310 | mem_ctrl_jal; // @[RocketCore.scala 747:35]
  assign io_imem_btb_update_bits_br_pc = _T_1776[38:0]; // @[RocketCore.scala 754:33]
  assign io_imem_btb_update_bits_cfiType = _T_1765 ? 2'h2 : _T_1772; // @[RocketCore.scala 748:35]
  assign io_imem_bht_update_valid = mem_reg_valid & ~take_pc_wb; // @[RocketCore.scala 758:28]
  assign io_imem_bht_update_bits_prediction_history = mem_reg_btb_resp_bht_history; // @[RocketCore.scala 763:38]
  assign io_imem_bht_update_bits_pc = io_imem_btb_update_bits_pc; // @[RocketCore.scala 759:30]
  assign io_imem_bht_update_bits_branch = mem_ctrl_branch; // @[RocketCore.scala 762:34]
  assign io_imem_bht_update_bits_taken = mem_br_taken; // @[RocketCore.scala 760:33]
  assign io_imem_bht_update_bits_mispredict = ex_pc_valid ? _T_1296 : _T_1299; // @[RocketCore.scala 761:38]
  assign io_imem_flush_icache = _T_1747 & ~io_dmem_s2_nack; // @[RocketCore.scala 732:24]
  assign io_dmem_req_valid = ex_reg_valid & ex_ctrl_mem; // @[RocketCore.scala 776:25]
  assign io_dmem_req_bits_addr = {msb_2,alu_io_adder_out[38:0]}; // @[RocketCore.scala 783:25]
  assign io_dmem_req_bits_tag = {{1'd0}, ex_dcache_tag}; // @[RocketCore.scala 779:25]
  assign io_dmem_req_bits_cmd = ex_ctrl_mem_cmd; // @[RocketCore.scala 780:25]
  assign io_dmem_req_bits_typ = ex_ctrl_mem_type; // @[RocketCore.scala 781:25]
  assign io_dmem_s1_kill = _T_1797 | fpu_kill_mem; // @[RocketCore.scala 785:19]
  assign io_dmem_s1_data_data = mem_ctrl_fp ? io_fpu_store_data : mem_reg_rs2; // @[RocketCore.scala 784:24]
  assign io_dmem_keep_clock_enabled = ibuf_io_inst_0_valid & id_ctrl_mem; // @[RocketCore.scala 788:30]
  assign io_ptw_ptbr_mode = csr_io_ptbr_mode; // @[RocketCore.scala 647:15]
  assign io_ptw_ptbr_ppn = csr_io_ptbr_ppn; // @[RocketCore.scala 647:15]
  assign io_ptw_sfence_valid = io_imem_sfence_valid; // @[RocketCore.scala 742:17]
  assign io_ptw_sfence_bits_rs1 = io_imem_sfence_bits_rs1; // @[RocketCore.scala 742:17]
  assign io_ptw_status_dprv = csr_io_status_dprv; // @[RocketCore.scala 649:17]
  assign io_ptw_status_prv = csr_io_status_prv; // @[RocketCore.scala 649:17]
  assign io_ptw_status_mxr = csr_io_status_mxr; // @[RocketCore.scala 649:17]
  assign io_ptw_status_sum = csr_io_status_sum; // @[RocketCore.scala 649:17]
  assign io_ptw_pmp_0_cfg_l = csr_io_pmp_0_cfg_l; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_0_cfg_a = csr_io_pmp_0_cfg_a; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_0_cfg_x = csr_io_pmp_0_cfg_x; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_0_cfg_w = csr_io_pmp_0_cfg_w; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_0_cfg_r = csr_io_pmp_0_cfg_r; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_0_addr = csr_io_pmp_0_addr; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_0_mask = csr_io_pmp_0_mask; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_1_cfg_l = csr_io_pmp_1_cfg_l; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_1_cfg_a = csr_io_pmp_1_cfg_a; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_1_cfg_x = csr_io_pmp_1_cfg_x; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_1_cfg_w = csr_io_pmp_1_cfg_w; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_1_cfg_r = csr_io_pmp_1_cfg_r; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_1_addr = csr_io_pmp_1_addr; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_1_mask = csr_io_pmp_1_mask; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_2_cfg_l = csr_io_pmp_2_cfg_l; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_2_cfg_a = csr_io_pmp_2_cfg_a; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_2_cfg_x = csr_io_pmp_2_cfg_x; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_2_cfg_w = csr_io_pmp_2_cfg_w; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_2_cfg_r = csr_io_pmp_2_cfg_r; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_2_addr = csr_io_pmp_2_addr; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_2_mask = csr_io_pmp_2_mask; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_3_cfg_l = csr_io_pmp_3_cfg_l; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_3_cfg_a = csr_io_pmp_3_cfg_a; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_3_cfg_x = csr_io_pmp_3_cfg_x; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_3_cfg_w = csr_io_pmp_3_cfg_w; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_3_cfg_r = csr_io_pmp_3_cfg_r; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_3_addr = csr_io_pmp_3_addr; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_3_mask = csr_io_pmp_3_mask; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_4_cfg_l = csr_io_pmp_4_cfg_l; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_4_cfg_a = csr_io_pmp_4_cfg_a; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_4_cfg_x = csr_io_pmp_4_cfg_x; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_4_cfg_w = csr_io_pmp_4_cfg_w; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_4_cfg_r = csr_io_pmp_4_cfg_r; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_4_addr = csr_io_pmp_4_addr; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_4_mask = csr_io_pmp_4_mask; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_5_cfg_l = csr_io_pmp_5_cfg_l; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_5_cfg_a = csr_io_pmp_5_cfg_a; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_5_cfg_x = csr_io_pmp_5_cfg_x; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_5_cfg_w = csr_io_pmp_5_cfg_w; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_5_cfg_r = csr_io_pmp_5_cfg_r; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_5_addr = csr_io_pmp_5_addr; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_5_mask = csr_io_pmp_5_mask; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_6_cfg_l = csr_io_pmp_6_cfg_l; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_6_cfg_a = csr_io_pmp_6_cfg_a; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_6_cfg_x = csr_io_pmp_6_cfg_x; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_6_cfg_w = csr_io_pmp_6_cfg_w; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_6_cfg_r = csr_io_pmp_6_cfg_r; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_6_addr = csr_io_pmp_6_addr; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_6_mask = csr_io_pmp_6_mask; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_7_cfg_l = csr_io_pmp_7_cfg_l; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_7_cfg_a = csr_io_pmp_7_cfg_a; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_7_cfg_x = csr_io_pmp_7_cfg_x; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_7_cfg_w = csr_io_pmp_7_cfg_w; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_7_cfg_r = csr_io_pmp_7_cfg_r; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_7_addr = csr_io_pmp_7_addr; // @[RocketCore.scala 650:14]
  assign io_ptw_pmp_7_mask = csr_io_pmp_7_mask; // @[RocketCore.scala 650:14]
  assign io_ptw_customCSRs_csrs_0_value = 64'h0; // @[RocketCore.scala 648:79]
  assign io_ptw_pcode_req_valid = csr_io_pcode_req_valid; // @[RocketCore.scala 268:20]
  assign io_ptw_pcode_req_bits_id = csr_io_pcode_req_bits_id; // @[RocketCore.scala 268:20]
  assign io_ptw_pcode_req_bits_value_base = csr_io_pcode_req_bits_value_base; // @[RocketCore.scala 268:20]
  assign io_ptw_pcode_req_bits_value_mask = csr_io_pcode_req_bits_value_mask; // @[RocketCore.scala 268:20]
  assign io_ptw_pcode_req_bits_value_valid = csr_io_pcode_req_bits_value_valid; // @[RocketCore.scala 268:20]
  assign io_ptw_pcode_req_bits_value_locked = csr_io_pcode_req_bits_value_locked; // @[RocketCore.scala 268:20]
  assign io_ptw_vpoffset_req_bits_value = csr_io_vpoffset_req_bits_value; // @[RocketCore.scala 271:23]
  assign io_fpu_inst = ibuf_io_inst_0_bits_inst_bits; // @[RocketCore.scala 768:15]
  assign io_fpu_fromint_data = ex_reg_rs_bypass_0 ? _T_981 : _T_982; // @[RocketCore.scala 769:23]
  assign io_fpu_fcsr_rm = csr_io_fcsr_rm; // @[RocketCore.scala 638:18]
  assign io_fpu_dmem_resp_val = dmem_resp_valid & io_dmem_resp_bits_tag[0]; // @[RocketCore.scala 770:24]
  assign io_fpu_dmem_resp_type = io_dmem_resp_bits_typ; // @[RocketCore.scala 772:25]
  assign io_fpu_dmem_resp_tag = io_dmem_resp_bits_tag[5:1]; // @[RocketCore.scala 773:24]
  assign io_fpu_dmem_resp_data = io_dmem_resp_bits_data_word_bypass; // @[RocketCore.scala 771:25]
  assign io_fpu_valid = ~ctrl_killd & id_ctrl_fp; // @[RocketCore.scala 765:16]
  assign io_fpu_killx = _T_1117 | ~ex_reg_valid; // @[RocketCore.scala 766:16]
  assign io_fpu_killm = _T_1418 | ~mem_reg_valid; // @[RocketCore.scala 767:16]
  assign ibuf_clock = clock;
  assign ibuf_reset = reset;
  assign ibuf_io_imem_valid = io_imem_resp_valid; // @[RocketCore.scala 240:16]
  assign ibuf_io_imem_bits_btb_taken = io_imem_resp_bits_btb_taken; // @[RocketCore.scala 240:16]
  assign ibuf_io_imem_bits_btb_bridx = io_imem_resp_bits_btb_bridx; // @[RocketCore.scala 240:16]
  assign ibuf_io_imem_bits_btb_entry = io_imem_resp_bits_btb_entry; // @[RocketCore.scala 240:16]
  assign ibuf_io_imem_bits_btb_bht_history = io_imem_resp_bits_btb_bht_history; // @[RocketCore.scala 240:16]
  assign ibuf_io_imem_bits_pc = io_imem_resp_bits_pc; // @[RocketCore.scala 240:16]
  assign ibuf_io_imem_bits_data = io_imem_resp_bits_data; // @[RocketCore.scala 240:16]
  assign ibuf_io_imem_bits_xcpt_pf_inst = io_imem_resp_bits_xcpt_pf_inst; // @[RocketCore.scala 240:16]
  assign ibuf_io_imem_bits_xcpt_ae_inst = io_imem_resp_bits_xcpt_ae_inst; // @[RocketCore.scala 240:16]
  assign ibuf_io_imem_bits_replay = io_imem_resp_bits_replay; // @[RocketCore.scala 240:16]
  assign ibuf_io_kill = take_pc_wb | take_pc_mem; // @[RocketCore.scala 241:16]
  assign ibuf_io_inst_0_ready = ~ctrl_stalld; // @[RocketCore.scala 744:25]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_ungated_clock = clock; // @[RocketCore.scala 630:24]
  assign csr_io_interrupts_debug = io_interrupts_debug; // @[RocketCore.scala 636:21]
  assign csr_io_interrupts_mtip = io_interrupts_mtip; // @[RocketCore.scala 636:21]
  assign csr_io_interrupts_msip = io_interrupts_msip; // @[RocketCore.scala 636:21]
  assign csr_io_interrupts_meip = io_interrupts_meip; // @[RocketCore.scala 636:21]
  assign csr_io_interrupts_seip = io_interrupts_seip; // @[RocketCore.scala 636:21]
  assign csr_io_hartid = io_hartid; // @[RocketCore.scala 637:17]
  assign csr_io_rw_addr = wb_reg_inst[31:20]; // @[RocketCore.scala 651:18]
  assign csr_io_rw_cmd = wb_ctrl_csr & ~_T_1540; // @[RocketCore.scala 652:17]
  assign csr_io_rw_wdata = wb_reg_wdata; // @[RocketCore.scala 653:19]
  assign csr_io_decode_0_csr = ibuf_io_inst_0_bits_raw[31:20]; // @[RocketCore.scala 631:24]
  assign csr_io_exception = _T_1453 | _T_1448; // @[RocketCore.scala 632:20]
  assign csr_io_retire = _T_1488 & ~wb_xcpt; // @[RocketCore.scala 634:17]
  assign csr_io_cause = wb_reg_xcpt ? wb_reg_cause : {{60'd0}, _T_1458}; // @[RocketCore.scala 633:16]
  assign csr_io_pc = wb_reg_pc; // @[RocketCore.scala 641:13]
  assign csr_io_tval = tval_valid ? _T_1537 : 40'h0; // @[RocketCore.scala 646:15]
  assign csr_io_fcsr_flags_valid = io_fpu_fcsr_flags_valid; // @[RocketCore.scala 639:21]
  assign csr_io_fcsr_flags_bits = io_fpu_fcsr_flags_bits; // @[RocketCore.scala 639:21]
  assign bpu_io_status_debug = csr_io_status_debug; // @[RocketCore.scala 303:17]
  assign bpu_io_status_prv = csr_io_status_prv; // @[RocketCore.scala 303:17]
  assign bpu_io_bp_0_control_action = csr_io_bp_0_control_action; // @[RocketCore.scala 304:13]
  assign bpu_io_bp_0_control_tmatch = csr_io_bp_0_control_tmatch; // @[RocketCore.scala 304:13]
  assign bpu_io_bp_0_control_m = csr_io_bp_0_control_m; // @[RocketCore.scala 304:13]
  assign bpu_io_bp_0_control_s = csr_io_bp_0_control_s; // @[RocketCore.scala 304:13]
  assign bpu_io_bp_0_control_u = csr_io_bp_0_control_u; // @[RocketCore.scala 304:13]
  assign bpu_io_bp_0_control_x = csr_io_bp_0_control_x; // @[RocketCore.scala 304:13]
  assign bpu_io_bp_0_control_w = csr_io_bp_0_control_w; // @[RocketCore.scala 304:13]
  assign bpu_io_bp_0_control_r = csr_io_bp_0_control_r; // @[RocketCore.scala 304:13]
  assign bpu_io_bp_0_address = csr_io_bp_0_address; // @[RocketCore.scala 304:13]
  assign bpu_io_pc = ibuf_io_pc[38:0]; // @[RocketCore.scala 305:13]
  assign bpu_io_ea = mem_reg_wdata[38:0]; // @[RocketCore.scala 306:13]
  assign alu_io_dw = ex_ctrl_alu_dw; // @[RocketCore.scala 362:13]
  assign alu_io_fn = ex_ctrl_alu_fn; // @[RocketCore.scala 363:13]
  assign alu_io_in2 = _T_1064 ? $signed(_T_1058) : $signed({{32{_T_1063[31]}},_T_1063}); // @[RocketCore.scala 364:14]
  assign alu_io_in1 = _T_1057 ? $signed(_T_1053) : $signed({{24{_T_1056[39]}},_T_1056}); // @[RocketCore.scala 365:14]
  assign div_clock = clock;
  assign div_reset = reset;
  assign div_io_req_valid = ex_reg_valid & ex_ctrl_div; // @[RocketCore.scala 377:20]
  assign div_io_req_bits_fn = ex_ctrl_alu_fn; // @[RocketCore.scala 379:22]
  assign div_io_req_bits_dw = ex_ctrl_alu_dw; // @[RocketCore.scala 378:22]
  assign div_io_req_bits_in1 = ex_reg_rs_bypass_0 ? _T_981 : _T_982; // @[RocketCore.scala 380:23]
  assign div_io_req_bits_in2 = ex_reg_rs_bypass_1 ? _T_989 : _T_990; // @[RocketCore.scala 381:23]
  assign div_io_req_bits_tag = ex_reg_inst[11:7]; // @[RocketCore.scala 382:23]
  assign div_io_kill = killm_common & _T_1422; // @[RocketCore.scala 541:15]
  assign div_io_resp_ready = _T_1486 ? 1'h0 : ~wb_wxd; // @[RocketCore.scala 597:21 RocketCore.scala 611:23]
  assign Rocket_cov_read_addr = Rocket_state;
  assign Rocket_cov_read_data = Rocket_cov[Rocket_cov_read_addr]; // @[Coverage map for Rocket]
  assign Rocket_cov_write_data = 1'h1;
  assign Rocket_cov_write_addr = Rocket_state;
  assign Rocket_cov_write_mask = 1'h1;
  assign Rocket_cov_write_en = 1'h1;
  assign mux_cond_0 = _T_1532;
  assign mux_cond_1 = _T_1501;
  assign mux_cond_2 = _T_1496;
  assign mux_cond_3 = _T_1500;
  assign mux_cond_4 = _T_1286;
  assign wb_ctrl_wfd_shl = {wb_ctrl_wfd, 1'h0};
  assign wb_ctrl_wfd_pad = {18'h0,wb_ctrl_wfd_shl};
  assign ex_ctrl_mem_type_shl = {ex_ctrl_mem_type, 4'h0};
  assign ex_ctrl_mem_type_pad = {13'h0,ex_ctrl_mem_type_shl};
  assign wb_reg_replay_shl = {wb_reg_replay, 8'h0};
  assign wb_reg_replay_pad = {11'h0,wb_reg_replay_shl};
  assign wb_ctrl_mem_shl = {wb_ctrl_mem, 19'h0};
  assign wb_ctrl_mem_pad = wb_ctrl_mem_shl;
  assign mem_ctrl_jalr_shl = {mem_ctrl_jalr, 11'h0};
  assign mem_ctrl_jalr_pad = {8'h0,mem_ctrl_jalr_shl};
  assign ex_ctrl_wfd_shl = {ex_ctrl_wfd, 3'h0};
  assign ex_ctrl_wfd_pad = {16'h0,ex_ctrl_wfd_shl};
  assign mem_ctrl_wfd_shl = {mem_ctrl_wfd, 1'h0};
  assign mem_ctrl_wfd_pad = {18'h0,mem_ctrl_wfd_shl};
  assign ex_ctrl_sel_alu1_shl = {ex_ctrl_sel_alu1, 14'h0};
  assign ex_ctrl_sel_alu1_pad = {4'h0,ex_ctrl_sel_alu1_shl};
  assign ex_ctrl_fp_shl = {ex_ctrl_fp, 19'h0};
  assign ex_ctrl_fp_pad = ex_ctrl_fp_shl;
  assign mem_reg_rvc_shl = {mem_reg_rvc, 2'h0};
  assign mem_reg_rvc_pad = {17'h0,mem_reg_rvc_shl};
  assign ex_ctrl_rxs2_shl = {ex_ctrl_rxs2, 5'h0};
  assign ex_ctrl_rxs2_pad = {14'h0,ex_ctrl_rxs2_shl};
  assign ex_reg_xcpt_interrupt_shl = {ex_reg_xcpt_interrupt, 3'h0};
  assign ex_reg_xcpt_interrupt_pad = {16'h0,ex_reg_xcpt_interrupt_shl};
  assign mem_reg_valid_shl = {mem_reg_valid, 4'h0};
  assign mem_reg_valid_pad = {15'h0,mem_reg_valid_shl};
  assign mem_ctrl_mem_shl = {mem_ctrl_mem, 6'h0};
  assign mem_ctrl_mem_pad = {13'h0,mem_ctrl_mem_shl};
  assign mem_reg_store_shl = mem_reg_store;
  assign mem_reg_store_pad = {19'h0,mem_reg_store_shl};
  assign mem_reg_xcpt_shl = {mem_reg_xcpt, 6'h0};
  assign mem_reg_xcpt_pad = {13'h0,mem_reg_xcpt_shl};
  assign mem_ctrl_branch_shl = {mem_ctrl_branch, 1'h0};
  assign mem_ctrl_branch_pad = {18'h0,mem_ctrl_branch_shl};
  assign ex_ctrl_wxd_shl = {ex_ctrl_wxd, 11'h0};
  assign ex_ctrl_wxd_pad = {8'h0,ex_ctrl_wxd_shl};
  assign mem_ctrl_wxd_shl = {mem_ctrl_wxd, 2'h0};
  assign mem_ctrl_wxd_pad = {17'h0,mem_ctrl_wxd_shl};
  assign ex_ctrl_mem_shl = {ex_ctrl_mem, 7'h0};
  assign ex_ctrl_mem_pad = {12'h0,ex_ctrl_mem_shl};
  assign mem_reg_replay_shl = {mem_reg_replay, 3'h0};
  assign mem_reg_replay_pad = {16'h0,mem_reg_replay_shl};
  assign wb_reg_xcpt_shl = {wb_reg_xcpt, 8'h0};
  assign wb_reg_xcpt_pad = {11'h0,wb_reg_xcpt_shl};
  assign mem_ctrl_jal_shl = {mem_ctrl_jal, 9'h0};
  assign mem_ctrl_jal_pad = {10'h0,mem_ctrl_jal_shl};
  assign ex_ctrl_jalr_shl = {ex_ctrl_jalr, 1'h0};
  assign ex_ctrl_jalr_pad = {18'h0,ex_ctrl_jalr_shl};
  assign mem_reg_flush_pipe_shl = {mem_reg_flush_pipe, 17'h0};
  assign mem_reg_flush_pipe_pad = {2'h0,mem_reg_flush_pipe_shl};
  assign mem_reg_xcpt_interrupt_shl = {mem_reg_xcpt_interrupt, 10'h0};
  assign mem_reg_xcpt_interrupt_pad = {9'h0,mem_reg_xcpt_interrupt_shl};
  assign ex_reg_replay_shl = {ex_reg_replay, 7'h0};
  assign ex_reg_replay_pad = {12'h0,ex_reg_replay_shl};
  assign ex_ctrl_sel_alu2_shl = {ex_ctrl_sel_alu2, 12'h0};
  assign ex_ctrl_sel_alu2_pad = {6'h0,ex_ctrl_sel_alu2_shl};
  assign ex_reg_valid_shl = {ex_reg_valid, 5'h0};
  assign ex_reg_valid_pad = {14'h0,ex_reg_valid_shl};
  assign mem_ctrl_fp_shl = {mem_ctrl_fp, 9'h0};
  assign mem_ctrl_fp_pad = {10'h0,mem_ctrl_fp_shl};
  assign id_reg_fence_shl = {id_reg_fence, 12'h0};
  assign id_reg_fence_pad = {7'h0,id_reg_fence_shl};
  assign wb_ctrl_div_shl = {wb_ctrl_div, 1'h0};
  assign wb_ctrl_div_pad = {18'h0,wb_ctrl_div_shl};
  assign ex_ctrl_sel_imm_shl = {ex_ctrl_sel_imm, 2'h0};
  assign ex_ctrl_sel_imm_pad = {15'h0,ex_ctrl_sel_imm_shl};
  assign wb_ctrl_wxd_shl = {wb_ctrl_wxd, 9'h0};
  assign wb_ctrl_wxd_pad = {10'h0,wb_ctrl_wxd_shl};
  assign ex_ctrl_div_shl = {ex_ctrl_div, 12'h0};
  assign ex_ctrl_div_pad = {7'h0,ex_ctrl_div_shl};
  assign wb_reg_valid_shl = {wb_reg_valid, 14'h0};
  assign wb_reg_valid_pad = {5'h0,wb_reg_valid_shl};
  assign mem_reg_sfence_shl = {mem_reg_sfence, 9'h0};
  assign mem_reg_sfence_pad = {10'h0,mem_reg_sfence_shl};
  assign ex_reg_rvc_shl = {ex_reg_rvc, 9'h0};
  assign ex_reg_rvc_pad = {10'h0,ex_reg_rvc_shl};
  assign mem_reg_load_shl = {mem_reg_load, 19'h0};
  assign mem_reg_load_pad = mem_reg_load_shl;
  assign wb_reg_flush_pipe_shl = {wb_reg_flush_pipe, 13'h0};
  assign wb_reg_flush_pipe_pad = {6'h0,wb_reg_flush_pipe_shl};
  assign mem_reg_slow_bypass_shl = {mem_reg_slow_bypass, 10'h0};
  assign mem_reg_slow_bypass_pad = {9'h0,mem_reg_slow_bypass_shl};
  assign blocked_shl = {blocked, 8'h0};
  assign blocked_pad = {11'h0,blocked_shl};
  assign mem_br_taken_shl = {mem_br_taken, 9'h0};
  assign mem_br_taken_pad = {10'h0,mem_br_taken_shl};
  assign mem_ctrl_div_shl = {mem_ctrl_div, 6'h0};
  assign mem_ctrl_div_pad = {13'h0,mem_ctrl_div_shl};
  assign mux_cond_0_shl = {mux_cond_0, 13'h0};
  assign mux_cond_0_pad = {6'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 15'h0};
  assign mux_cond_1_pad = {4'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 7'h0};
  assign mux_cond_2_pad = {12'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 8'h0};
  assign mux_cond_3_pad = {11'h0,mux_cond_3_shl};
  assign mux_cond_4_shl = {mux_cond_4, 1'h0};
  assign mux_cond_4_pad = {18'h0,mux_cond_4_shl};
  assign ex_reg_rs_bypass_0_shl = {ex_reg_rs_bypass_0, 8'h0};
  assign ex_reg_rs_bypass_0_pad = {11'h0,ex_reg_rs_bypass_0_shl};
  assign ex_reg_rs_bypass_1_shl = {ex_reg_rs_bypass_1, 8'h0};
  assign ex_reg_rs_bypass_1_pad = {11'h0,ex_reg_rs_bypass_1_shl};
  assign ex_reg_rs_lsb_0_shl = {ex_reg_rs_lsb_0, 17'h0};
  assign ex_reg_rs_lsb_0_pad = {1'h0,ex_reg_rs_lsb_0_shl};
  assign ex_reg_rs_lsb_1_shl = {ex_reg_rs_lsb_1, 17'h0};
  assign ex_reg_rs_lsb_1_pad = {1'h0,ex_reg_rs_lsb_1_shl};
  assign Rocket_xor32 = ex_ctrl_mem_type_pad ^ wb_reg_replay_pad;
  assign Rocket_xor15 = wb_ctrl_wfd_pad ^ Rocket_xor32;
  assign Rocket_xor34 = mem_ctrl_jalr_pad ^ ex_ctrl_wfd_pad;
  assign Rocket_xor16 = wb_ctrl_mem_pad ^ Rocket_xor34;
  assign Rocket_xor7 = Rocket_xor15 ^ Rocket_xor16;
  assign Rocket_xor36 = ex_ctrl_sel_alu1_pad ^ ex_ctrl_fp_pad;
  assign Rocket_xor17 = mem_ctrl_wfd_pad ^ Rocket_xor36;
  assign Rocket_xor37 = mem_reg_rvc_pad ^ ex_ctrl_rxs2_pad;
  assign Rocket_xor38 = ex_reg_xcpt_interrupt_pad ^ mem_reg_valid_pad;
  assign Rocket_xor18 = Rocket_xor37 ^ Rocket_xor38;
  assign Rocket_xor8 = Rocket_xor17 ^ Rocket_xor18;
  assign Rocket_xor3 = Rocket_xor7 ^ Rocket_xor8;
  assign Rocket_xor40 = mem_reg_store_pad ^ mem_reg_xcpt_pad;
  assign Rocket_xor19 = mem_ctrl_mem_pad ^ Rocket_xor40;
  assign Rocket_xor42 = ex_ctrl_wxd_pad ^ mem_ctrl_wxd_pad;
  assign Rocket_xor20 = mem_ctrl_branch_pad ^ Rocket_xor42;
  assign Rocket_xor9 = Rocket_xor19 ^ Rocket_xor20;
  assign Rocket_xor44 = mem_reg_replay_pad ^ wb_reg_xcpt_pad;
  assign Rocket_xor21 = ex_ctrl_mem_pad ^ Rocket_xor44;
  assign Rocket_xor45 = mem_ctrl_jal_pad ^ ex_ctrl_jalr_pad;
  assign Rocket_xor46 = mem_reg_flush_pipe_pad ^ mem_reg_xcpt_interrupt_pad;
  assign Rocket_xor22 = Rocket_xor45 ^ Rocket_xor46;
  assign Rocket_xor10 = Rocket_xor21 ^ Rocket_xor22;
  assign Rocket_xor4 = Rocket_xor9 ^ Rocket_xor10;
  assign Rocket_xor1 = Rocket_xor3 ^ Rocket_xor4;
  assign Rocket_xor48 = ex_ctrl_sel_alu2_pad ^ ex_reg_valid_pad;
  assign Rocket_xor23 = ex_reg_replay_pad ^ Rocket_xor48;
  assign Rocket_xor50 = id_reg_fence_pad ^ wb_ctrl_div_pad;
  assign Rocket_xor24 = mem_ctrl_fp_pad ^ Rocket_xor50;
  assign Rocket_xor11 = Rocket_xor23 ^ Rocket_xor24;
  assign Rocket_xor52 = wb_ctrl_wxd_pad ^ ex_ctrl_div_pad;
  assign Rocket_xor25 = ex_ctrl_sel_imm_pad ^ Rocket_xor52;
  assign Rocket_xor53 = wb_reg_valid_pad ^ mem_reg_sfence_pad;
  assign Rocket_xor54 = ex_reg_rvc_pad ^ mem_reg_load_pad;
  assign Rocket_xor26 = Rocket_xor53 ^ Rocket_xor54;
  assign Rocket_xor12 = Rocket_xor25 ^ Rocket_xor26;
  assign Rocket_xor5 = Rocket_xor11 ^ Rocket_xor12;
  assign Rocket_xor56 = mem_reg_slow_bypass_pad ^ blocked_pad;
  assign Rocket_xor27 = wb_reg_flush_pipe_pad ^ Rocket_xor56;
  assign Rocket_xor57 = mem_br_taken_pad ^ mem_ctrl_div_pad;
  assign Rocket_xor58 = mux_cond_0_pad ^ mux_cond_1_pad;
  assign Rocket_xor28 = Rocket_xor57 ^ Rocket_xor58;
  assign Rocket_xor13 = Rocket_xor27 ^ Rocket_xor28;
  assign Rocket_xor60 = mux_cond_3_pad ^ mux_cond_4_pad;
  assign Rocket_xor29 = mux_cond_2_pad ^ Rocket_xor60;
  assign Rocket_xor61 = ex_reg_rs_bypass_0_pad ^ ex_reg_rs_bypass_1_pad;
  assign Rocket_xor62 = ex_reg_rs_lsb_0_pad ^ ex_reg_rs_lsb_1_pad;
  assign Rocket_xor30 = Rocket_xor61 ^ Rocket_xor62;
  assign Rocket_xor14 = Rocket_xor29 ^ Rocket_xor30;
  assign Rocket_xor6 = Rocket_xor13 ^ Rocket_xor14;
  assign Rocket_xor2 = Rocket_xor5 ^ Rocket_xor6;
  assign Rocket_xor0 = Rocket_xor1 ^ Rocket_xor2;
  assign csr_sum = Rocket_covSum + csr_io_covSum;
  assign div_sum = csr_sum + div_io_covSum;
  assign ibuf_sum = div_sum + ibuf_io_covSum;
  assign alu_sum = ibuf_sum + alu_io_covSum;
  assign bpu_sum = alu_sum + bpu_io_covSum;
  assign io_covSum = bpu_sum;
  assign alu_metaAssert_wire = alu_metaAssert;
  assign bpu_metaAssert_wire = bpu_metaAssert;
  assign ibuf_metaAssert_wire = ibuf_metaAssert;
  assign csr_metaAssert_wire = csr_metaAssert;
  assign div_metaAssert_wire = div_metaAssert;
  assign Rocket_or1 = ibuf_metaAssert_wire | alu_metaAssert_wire;
  assign Rocket_or6 = div_metaAssert_wire | csr_metaAssert_wire;
  assign Rocket_or2 = bpu_metaAssert_wire | Rocket_or6;
  assign Rocket_or0 = Rocket_or1 | Rocket_or2;
  assign metaAssert = Rocket_metaAssert;
  assign csr_metaReset = metaReset | csr_halt;
  assign div_metaReset = metaReset | div_halt;
  assign ibuf_metaReset = metaReset | ibuf_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 31; initvar = initvar+1)
    _T_760[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{`RANDOM}};
  _RAND_2 = {2{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  imem_might_request_reg = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  ex_ctrl_fp = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  ex_ctrl_branch = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  ex_ctrl_jal = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ex_ctrl_jalr = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  ex_ctrl_rxs2 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  ex_ctrl_sel_alu2 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  ex_ctrl_sel_alu1 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  ex_ctrl_sel_imm = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  ex_ctrl_alu_dw = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  ex_ctrl_alu_fn = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  ex_ctrl_mem = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  ex_ctrl_mem_cmd = _RAND_15[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  ex_ctrl_mem_type = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  ex_ctrl_wfd = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  ex_ctrl_div = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  ex_ctrl_wxd = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  ex_ctrl_csr = _RAND_20[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  ex_ctrl_fence_i = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  mem_ctrl_fp = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  mem_ctrl_branch = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  mem_ctrl_jal = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  mem_ctrl_jalr = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  mem_ctrl_mem = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  mem_ctrl_mem_type = _RAND_27[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  mem_ctrl_wfd = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  mem_ctrl_div = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  mem_ctrl_wxd = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  mem_ctrl_csr = _RAND_31[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  mem_ctrl_fence_i = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  wb_ctrl_mem = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  wb_ctrl_mem_type = _RAND_34[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  wb_ctrl_wfd = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  wb_ctrl_div = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  wb_ctrl_wxd = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  wb_ctrl_csr = _RAND_38[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  wb_ctrl_fence_i = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  ex_reg_xcpt_interrupt = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  ex_reg_valid = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  ex_reg_rvc = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  ex_reg_btb_resp_entry = _RAND_43[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  ex_reg_btb_resp_bht_history = _RAND_44[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  ex_reg_xcpt = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  ex_reg_flush_pipe = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  ex_reg_load_use = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {2{`RANDOM}};
  ex_reg_cause = _RAND_48[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  ex_reg_replay = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {2{`RANDOM}};
  ex_reg_pc = _RAND_50[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  ex_reg_inst = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  mem_reg_xcpt_interrupt = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  mem_reg_valid = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  mem_reg_rvc = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  mem_reg_btb_resp_entry = _RAND_55[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  mem_reg_btb_resp_bht_history = _RAND_56[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  mem_reg_xcpt = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  mem_reg_replay = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  mem_reg_flush_pipe = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {2{`RANDOM}};
  mem_reg_cause = _RAND_60[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  mem_reg_slow_bypass = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  mem_reg_load = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  mem_reg_store = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  mem_reg_sfence = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {2{`RANDOM}};
  mem_reg_pc = _RAND_65[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  mem_reg_inst = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {2{`RANDOM}};
  mem_reg_wdata = _RAND_67[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {2{`RANDOM}};
  mem_reg_rs2 = _RAND_68[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  mem_br_taken = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  wb_reg_valid = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  wb_reg_xcpt = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  wb_reg_replay = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  wb_reg_flush_pipe = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {2{`RANDOM}};
  wb_reg_cause = _RAND_74[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  wb_reg_sfence = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {2{`RANDOM}};
  wb_reg_pc = _RAND_76[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  wb_reg_inst = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {2{`RANDOM}};
  wb_reg_wdata = _RAND_78[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  id_reg_fence = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  ex_reg_rs_bypass_0 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  ex_reg_rs_bypass_1 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  ex_reg_rs_lsb_0 = _RAND_82[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  ex_reg_rs_lsb_1 = _RAND_83[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {2{`RANDOM}};
  ex_reg_rs_msb_0 = _RAND_84[61:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {2{`RANDOM}};
  ex_reg_rs_msb_1 = _RAND_85[61:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_1550 = _RAND_86[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_1663 = _RAND_87[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  blocked = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_1422 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  Rocket_state = _RAND_90[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    Rocket_cov[initvar] = _RAND_91[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  Rocket_covSum = _RAND_92[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  Rocket_metaAssert = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_760__T_1499_en & _T_760__T_1499_mask) begin
      _T_760[_T_760__T_1499_addr] <= _T_760__T_1499_data; // @[RocketCore.scala 932:23]
    end
    if (metaReset) begin
      imem_might_request_reg <= 1'h0;
    end else begin
      imem_might_request_reg <= _T_1750 | io_ptw_customCSRs_csrs_0_value[1];
    end
    if (metaReset) begin
      ex_ctrl_fp <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_fp <= id_ctrl_fp;
    end
    if (metaReset) begin
      ex_ctrl_branch <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_branch <= id_ctrl_branch;
    end
    if (metaReset) begin
      ex_ctrl_jal <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_jal <= id_ctrl_jal;
    end
    if (metaReset) begin
      ex_ctrl_jalr <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_jalr <= id_ctrl_jalr;
    end
    if (metaReset) begin
      ex_ctrl_rxs2 <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_rxs2 <= id_ctrl_rxs2;
    end
    if (metaReset) begin
      ex_ctrl_sel_alu2 <= 2'h0;
    end else if (~ctrl_killd) begin
      if (id_xcpt) begin
        if (_T_1082) begin
          ex_ctrl_sel_alu2 <= 2'h0;
        end else if (_T_1079) begin
          ex_ctrl_sel_alu2 <= 2'h1;
        end else begin
          ex_ctrl_sel_alu2 <= 2'h0;
        end
      end else begin
        ex_ctrl_sel_alu2 <= id_ctrl_sel_alu2;
      end
    end
    if (metaReset) begin
      ex_ctrl_sel_alu1 <= 2'h0;
    end else if (~ctrl_killd) begin
      if (id_xcpt) begin
        if (_T_1082) begin
          ex_ctrl_sel_alu1 <= 2'h2;
        end else if (_T_1079) begin
          ex_ctrl_sel_alu1 <= 2'h2;
        end else begin
          ex_ctrl_sel_alu1 <= 2'h1;
        end
      end else begin
        ex_ctrl_sel_alu1 <= id_ctrl_sel_alu1;
      end
    end
    if (metaReset) begin
      ex_ctrl_sel_imm <= 3'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_sel_imm <= id_ctrl_sel_imm;
    end
    if (metaReset) begin
      ex_ctrl_alu_dw <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_alu_dw <= _GEN_8;
    end
    if (metaReset) begin
      ex_ctrl_alu_fn <= 4'h0;
    end else if (~ctrl_killd) begin
      if (id_xcpt) begin
        ex_ctrl_alu_fn <= 4'h0;
      end else begin
        ex_ctrl_alu_fn <= id_ctrl_alu_fn;
      end
    end
    if (metaReset) begin
      ex_ctrl_mem <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_mem <= id_ctrl_mem;
    end
    if (metaReset) begin
      ex_ctrl_mem_cmd <= 5'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_mem_cmd <= id_ctrl_mem_cmd;
    end
    if (metaReset) begin
      ex_ctrl_mem_type <= 3'h0;
    end else if (~ctrl_killd) begin
      if (id_sfence) begin
        ex_ctrl_mem_type <= {{1'd0}, _T_1086};
      end else begin
        ex_ctrl_mem_type <= id_ctrl_mem_type;
      end
    end
    if (metaReset) begin
      ex_ctrl_wfd <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_wfd <= id_ctrl_wfd;
    end
    if (metaReset) begin
      ex_ctrl_div <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_div <= id_ctrl_div;
    end
    if (metaReset) begin
      ex_ctrl_wxd <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_wxd <= id_ctrl_wxd;
    end
    if (metaReset) begin
      ex_ctrl_csr <= 3'h0;
    end else if (~ctrl_killd) begin
      if (id_csr_ren) begin
        ex_ctrl_csr <= 3'h2;
      end else begin
        ex_ctrl_csr <= id_ctrl_csr;
      end
    end
    if (metaReset) begin
      ex_ctrl_fence_i <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_fence_i <= id_ctrl_fence_i;
    end
    if (metaReset) begin
      mem_ctrl_fp <= 1'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_ctrl_fp <= ex_ctrl_fp;
      end
    end
    if (metaReset) begin
      mem_ctrl_branch <= 1'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_ctrl_branch <= ex_ctrl_branch;
      end
    end
    if (metaReset) begin
      mem_ctrl_jal <= 1'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_ctrl_jal <= ex_ctrl_jal;
      end
    end
    if (metaReset) begin
      mem_ctrl_jalr <= 1'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_ctrl_jalr <= ex_ctrl_jalr;
      end
    end
    if (metaReset) begin
      mem_ctrl_mem <= 1'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_ctrl_mem <= ex_ctrl_mem;
      end
    end
    if (metaReset) begin
      mem_ctrl_mem_type <= 3'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_ctrl_mem_type <= ex_ctrl_mem_type;
      end
    end
    if (metaReset) begin
      mem_ctrl_wfd <= 1'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_ctrl_wfd <= ex_ctrl_wfd;
      end
    end
    if (metaReset) begin
      mem_ctrl_div <= 1'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_ctrl_div <= ex_ctrl_div;
      end
    end
    if (metaReset) begin
      mem_ctrl_wxd <= 1'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_ctrl_wxd <= ex_ctrl_wxd;
      end
    end
    if (metaReset) begin
      mem_ctrl_csr <= 3'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_ctrl_csr <= ex_ctrl_csr;
      end
    end
    if (metaReset) begin
      mem_ctrl_fence_i <= 1'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_ctrl_fence_i <= _GEN_72;
      end
    end
    if (metaReset) begin
      wb_ctrl_mem <= 1'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_mem <= mem_ctrl_mem;
    end
    if (metaReset) begin
      wb_ctrl_mem_type <= 3'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_mem_type <= mem_ctrl_mem_type;
    end
    if (metaReset) begin
      wb_ctrl_wfd <= 1'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_wfd <= mem_ctrl_wfd;
    end
    if (metaReset) begin
      wb_ctrl_div <= 1'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_div <= mem_ctrl_div;
    end
    if (metaReset) begin
      wb_ctrl_wxd <= 1'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_wxd <= mem_ctrl_wxd;
    end
    if (metaReset) begin
      wb_ctrl_csr <= 3'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_csr <= mem_ctrl_csr;
    end
    if (metaReset) begin
      wb_ctrl_fence_i <= 1'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_fence_i <= mem_ctrl_fence_i;
    end
    if (metaReset) begin
      ex_reg_xcpt_interrupt <= 1'h0;
    end else begin
      ex_reg_xcpt_interrupt <= _T_1070 & csr_io_interrupt;
    end
    if (metaReset) begin
      ex_reg_valid <= 1'h0;
    end else begin
      ex_reg_valid <= ~ctrl_killd;
    end
    if (metaReset) begin
      ex_reg_rvc <= 1'h0;
    end else if (~ctrl_killd) begin
      if (id_xcpt) begin
        ex_reg_rvc <= _GEN_4;
      end else begin
        ex_reg_rvc <= ibuf_io_inst_0_bits_rvc;
      end
    end
    if (metaReset) begin
      ex_reg_btb_resp_entry <= 5'h0;
    end else if (_T_1108) begin
      ex_reg_btb_resp_entry <= ibuf_io_btb_resp_entry;
    end
    if (metaReset) begin
      ex_reg_btb_resp_bht_history <= 8'h0;
    end else if (_T_1108) begin
      ex_reg_btb_resp_bht_history <= ibuf_io_btb_resp_bht_history;
    end
    if (metaReset) begin
      ex_reg_xcpt <= 1'h0;
    end else begin
      ex_reg_xcpt <= ~ctrl_killd & id_xcpt;
    end
    if (metaReset) begin
      ex_reg_flush_pipe <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_reg_flush_pipe <= _T_1083;
    end
    if (metaReset) begin
      ex_reg_load_use <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_reg_load_use <= id_load_use;
    end
    if (metaReset) begin
      ex_reg_cause <= 64'h0;
    end else if (_T_1108) begin
      if (csr_io_interrupt) begin
        ex_reg_cause <= csr_io_interrupt_cause;
      end else begin
        ex_reg_cause <= {{60'd0}, _T_923};
      end
    end
    if (metaReset) begin
      ex_reg_replay <= 1'h0;
    end else begin
      ex_reg_replay <= _T_1070 & ibuf_io_inst_0_bits_replay;
    end
    if (metaReset) begin
      ex_reg_pc <= 40'h0;
    end else if (_T_1108) begin
      ex_reg_pc <= ibuf_io_pc;
    end
    if (metaReset) begin
      ex_reg_inst <= 32'h0;
    end else if (_T_1108) begin
      ex_reg_inst <= ibuf_io_inst_0_bits_inst_bits;
    end
    if (metaReset) begin
      mem_reg_xcpt_interrupt <= 1'h0;
    end else begin
      mem_reg_xcpt_interrupt <= ~take_pc_mem_wb & ex_reg_xcpt_interrupt;
    end
    if (metaReset) begin
      mem_reg_valid <= 1'h0;
    end else begin
      mem_reg_valid <= ~ctrl_killx;
    end
    if (metaReset) begin
      mem_reg_rvc <= 1'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_reg_rvc <= ex_reg_rvc;
      end
    end
    if (metaReset) begin
      mem_reg_btb_resp_entry <= 5'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_reg_btb_resp_entry <= ex_reg_btb_resp_entry;
      end
    end
    if (metaReset) begin
      mem_reg_btb_resp_bht_history <= 8'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_reg_btb_resp_bht_history <= ex_reg_btb_resp_bht_history;
      end
    end
    if (metaReset) begin
      mem_reg_xcpt <= 1'h0;
    end else begin
      mem_reg_xcpt <= ~ctrl_killx & ex_xcpt;
    end
    if (metaReset) begin
      mem_reg_replay <= 1'h0;
    end else begin
      mem_reg_replay <= ~take_pc_mem_wb & replay_ex;
    end
    if (metaReset) begin
      mem_reg_flush_pipe <= 1'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_reg_flush_pipe <= _GEN_73;
      end
    end
    if (metaReset) begin
      mem_reg_cause <= 64'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_reg_cause <= ex_reg_cause;
      end
    end
    if (metaReset) begin
      mem_reg_slow_bypass <= 1'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_reg_slow_bypass <= ex_slow_bypass;
      end
    end
    if (metaReset) begin
      mem_reg_load <= 1'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_reg_load <= _T_1348;
      end
    end
    if (metaReset) begin
      mem_reg_store <= 1'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_reg_store <= _T_1372;
      end
    end
    if (metaReset) begin
      mem_reg_sfence <= 1'h0;
    end else if (_T_1324) begin
      mem_reg_sfence <= 1'h0;
    end else if (ex_pc_valid) begin
      mem_reg_sfence <= ex_sfence;
    end
    if (metaReset) begin
      mem_reg_pc <= 40'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_reg_pc <= ex_reg_pc;
      end
    end
    if (metaReset) begin
      mem_reg_inst <= 32'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_reg_inst <= ex_reg_inst;
      end
    end
    if (metaReset) begin
      mem_reg_wdata <= 64'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_reg_wdata <= alu_io_out;
      end
    end
    if (metaReset) begin
      mem_reg_rs2 <= 64'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        if (_T_1375) begin
          if (_T_1377) begin
            mem_reg_rs2 <= _T_1381;
          end else if (_T_1382) begin
            mem_reg_rs2 <= _T_1385;
          end else if (_T_1386) begin
            mem_reg_rs2 <= _T_1388;
          end else if (ex_reg_rs_bypass_1) begin
            if (_T_988) begin
              mem_reg_rs2 <= io_dmem_resp_bits_data_word_bypass;
            end else if (_T_986) begin
              mem_reg_rs2 <= wb_reg_wdata;
            end else if (_T_984) begin
              mem_reg_rs2 <= mem_reg_wdata;
            end else begin
              mem_reg_rs2 <= 64'h0;
            end
          end else begin
            mem_reg_rs2 <= _T_990;
          end
        end
      end
    end
    if (metaReset) begin
      mem_br_taken <= 1'h0;
    end else if (!(_T_1324)) begin
      if (ex_pc_valid) begin
        mem_br_taken <= alu_io_cmp_out;
      end
    end
    if (metaReset) begin
      wb_reg_valid <= 1'h0;
    end else begin
      wb_reg_valid <= ~ctrl_killm;
    end
    if (metaReset) begin
      wb_reg_xcpt <= 1'h0;
    end else begin
      wb_reg_xcpt <= mem_xcpt & ~take_pc_wb;
    end
    if (metaReset) begin
      wb_reg_replay <= 1'h0;
    end else begin
      wb_reg_replay <= replay_mem & ~take_pc_wb;
    end
    if (metaReset) begin
      wb_reg_flush_pipe <= 1'h0;
    end else begin
      wb_reg_flush_pipe <= ~ctrl_killm & mem_reg_flush_pipe;
    end
    if (metaReset) begin
      wb_reg_cause <= 64'h0;
    end else if (mem_pc_valid) begin
      if (_T_1397) begin
        wb_reg_cause <= mem_reg_cause;
      end else begin
        wb_reg_cause <= {{60'd0}, _T_1401};
      end
    end
    if (metaReset) begin
      wb_reg_sfence <= 1'h0;
    end else if (mem_pc_valid) begin
      wb_reg_sfence <= mem_reg_sfence;
    end
    if (metaReset) begin
      wb_reg_pc <= 40'h0;
    end else if (mem_pc_valid) begin
      wb_reg_pc <= mem_reg_pc;
    end
    if (metaReset) begin
      wb_reg_inst <= 32'h0;
    end else if (mem_pc_valid) begin
      wb_reg_inst <= mem_reg_inst;
    end
    if (metaReset) begin
      wb_reg_wdata <= 64'h0;
    end else if (mem_pc_valid) begin
      if (_T_1434) begin
        wb_reg_wdata <= io_fpu_toint_data;
      end else begin
        wb_reg_wdata <= mem_int_wdata;
      end
    end
    if (metaReset) begin
      id_reg_fence <= 1'h0;
    end else if (reset) begin
      id_reg_fence <= 1'h0;
    end else if (~ctrl_killd) begin
      id_reg_fence <= _GEN_1;
    end else if (~id_mem_busy) begin
      id_reg_fence <= 1'h0;
    end
    if (metaReset) begin
      ex_reg_rs_bypass_0 <= 1'h0;
    end else if (~ctrl_killd) begin
      if (id_illegal_insn) begin
        ex_reg_rs_bypass_0 <= 1'h0;
      end else begin
        ex_reg_rs_bypass_0 <= do_bypass;
      end
    end
    if (metaReset) begin
      ex_reg_rs_bypass_1 <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_reg_rs_bypass_1 <= do_bypass_1;
    end
    if (metaReset) begin
      ex_reg_rs_lsb_0 <= 2'h0;
    end else if (~ctrl_killd) begin
      if (id_illegal_insn) begin
        ex_reg_rs_lsb_0 <= inst[1:0];
      end else if (_T_1092) begin
        ex_reg_rs_lsb_0 <= _GEN_228[1:0];
      end else if (_T_939) begin
        ex_reg_rs_lsb_0 <= 2'h0;
      end else if (_T_942) begin
        ex_reg_rs_lsb_0 <= 2'h1;
      end else if (_T_944) begin
        ex_reg_rs_lsb_0 <= 2'h2;
      end else begin
        ex_reg_rs_lsb_0 <= 2'h3;
      end
    end
    if (metaReset) begin
      ex_reg_rs_lsb_1 <= 2'h0;
    end else if (~ctrl_killd) begin
      if (_T_1100) begin
        ex_reg_rs_lsb_1 <= _GEN_229[1:0];
      end else if (_T_947) begin
        ex_reg_rs_lsb_1 <= 2'h0;
      end else if (_T_950) begin
        ex_reg_rs_lsb_1 <= 2'h1;
      end else if (_T_952) begin
        ex_reg_rs_lsb_1 <= 2'h2;
      end else begin
        ex_reg_rs_lsb_1 <= 2'h3;
      end
    end
    if (metaReset) begin
      ex_reg_rs_msb_0 <= 62'h0;
    end else if (~ctrl_killd) begin
      if (id_illegal_insn) begin
        ex_reg_rs_msb_0 <= {{32'd0}, inst[31:2]};
      end else if (_T_1092) begin
        ex_reg_rs_msb_0 <= _GEN_228[63:2];
      end
    end
    if (metaReset) begin
      ex_reg_rs_msb_1 <= 62'h0;
    end else if (~ctrl_killd) begin
      if (_T_1100) begin
        ex_reg_rs_msb_1 <= _GEN_229[63:2];
      end
    end
    if (metaReset) begin
      _T_1550 <= 32'h0;
    end else if (reset) begin
      _T_1550 <= 32'h0;
    end else if (_T_1584) begin
      _T_1550 <= _T_1583;
    end else if (ll_wen) begin
      _T_1550 <= _T_1556;
    end
    if (metaReset) begin
      _T_1663 <= 32'h0;
    end else if (reset) begin
      _T_1663 <= 32'h0;
    end else if (_T_1681) begin
      _T_1663 <= _T_1680;
    end else if (_T_1676) begin
      _T_1663 <= _T_1675;
    end else if (_T_1666) begin
      _T_1663 <= _T_1669;
    end
    if (metaReset) begin
      blocked <= 1'h0;
    end else begin
      blocked <= _T_1700 & _T_1702;
    end
    if (metaReset) begin
      _T_1422 <= 1'h0;
    end else begin
      _T_1422 <= div_io_req_ready & div_io_req_valid;
    end
    Rocket_state <= Rocket_xor0;
    if (!(Rocket_cov_read_data)) begin
      Rocket_covSum <= Rocket_covSum + 1'h1;
    end
    if (metaReset) begin
      Rocket_metaAssert <= 1'h0;
    end else begin
      Rocket_metaAssert <= Rocket_metaAssert | Rocket_or0;
    end
  end
  always @(posedge clock) begin
    if(Rocket_cov_write_en & Rocket_cov_write_mask) begin
      Rocket_cov[Rocket_cov_write_addr] <= Rocket_cov_write_data; // @[Coverage map for Rocket]
    end
  end
endmodule
module TLMonitor_64(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_param,
  input  [3:0]  io_in_a_bits_size,
  input         io_in_a_bits_source,
  input  [31:0] io_in_a_bits_address,
  input  [7:0]  io_in_a_bits_mask,
  input         io_in_b_ready,
  input         io_in_b_valid,
  input  [2:0]  io_in_b_bits_opcode,
  input  [1:0]  io_in_b_bits_param,
  input  [3:0]  io_in_b_bits_size,
  input         io_in_b_bits_source,
  input  [31:0] io_in_b_bits_address,
  input  [7:0]  io_in_b_bits_mask,
  input         io_in_b_bits_corrupt,
  input         io_in_c_ready,
  input         io_in_c_valid,
  input  [2:0]  io_in_c_bits_opcode,
  input  [2:0]  io_in_c_bits_param,
  input  [3:0]  io_in_c_bits_size,
  input         io_in_c_bits_source,
  input  [31:0] io_in_c_bits_address,
  input         io_in_d_ready,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [1:0]  io_in_d_bits_param,
  input  [3:0]  io_in_d_bits_size,
  input         io_in_d_bits_source,
  input  [1:0]  io_in_d_bits_sink,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt,
  input         io_in_e_ready,
  input         io_in_e_valid,
  input  [1:0]  io_in_e_bits_sink,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire  _T_30; // @[Parameters.scala 280:46]
  wire [26:0] _T_32; // @[package.scala 185:77]
  wire [31:0] _GEN_33; // @[Edges.scala 21:16]
  wire [31:0] _T_35; // @[Edges.scala 21:16]
  wire  _T_36; // @[Edges.scala 21:24]
  wire [3:0] _T_39; // @[OneHot.scala 52:12]
  wire [2:0] _T_41; // @[Misc.scala 206:81]
  wire  _T_42; // @[Misc.scala 210:21]
  wire  _T_47; // @[Misc.scala 219:38]
  wire  _T_48; // @[Misc.scala 219:29]
  wire  _T_50; // @[Misc.scala 219:38]
  wire  _T_51; // @[Misc.scala 219:29]
  wire  _T_55; // @[Misc.scala 218:27]
  wire  _T_56; // @[Misc.scala 219:38]
  wire  _T_57; // @[Misc.scala 219:29]
  wire  _T_58; // @[Misc.scala 218:27]
  wire  _T_59; // @[Misc.scala 219:38]
  wire  _T_60; // @[Misc.scala 219:29]
  wire  _T_61; // @[Misc.scala 218:27]
  wire  _T_62; // @[Misc.scala 219:38]
  wire  _T_63; // @[Misc.scala 219:29]
  wire  _T_64; // @[Misc.scala 218:27]
  wire  _T_65; // @[Misc.scala 219:38]
  wire  _T_66; // @[Misc.scala 219:29]
  wire  _T_70; // @[Misc.scala 218:27]
  wire  _T_71; // @[Misc.scala 219:38]
  wire  _T_72; // @[Misc.scala 219:29]
  wire  _T_73; // @[Misc.scala 218:27]
  wire  _T_74; // @[Misc.scala 219:38]
  wire  _T_75; // @[Misc.scala 219:29]
  wire  _T_76; // @[Misc.scala 218:27]
  wire  _T_77; // @[Misc.scala 219:38]
  wire  _T_78; // @[Misc.scala 219:29]
  wire  _T_79; // @[Misc.scala 218:27]
  wire  _T_80; // @[Misc.scala 219:38]
  wire  _T_81; // @[Misc.scala 219:29]
  wire  _T_82; // @[Misc.scala 218:27]
  wire  _T_83; // @[Misc.scala 219:38]
  wire  _T_84; // @[Misc.scala 219:29]
  wire  _T_85; // @[Misc.scala 218:27]
  wire  _T_86; // @[Misc.scala 219:38]
  wire  _T_87; // @[Misc.scala 219:29]
  wire  _T_88; // @[Misc.scala 218:27]
  wire  _T_89; // @[Misc.scala 219:38]
  wire  _T_90; // @[Misc.scala 219:29]
  wire  _T_91; // @[Misc.scala 218:27]
  wire  _T_92; // @[Misc.scala 219:38]
  wire  _T_93; // @[Misc.scala 219:29]
  wire [7:0] _T_100; // @[Cat.scala 30:58]
  wire [32:0] _T_104; // @[Parameters.scala 121:49]
  wire  _T_121; // @[Monitor.scala 48:25]
  wire  _T_123; // @[Parameters.scala 90:42]
  wire [31:0] _T_126; // @[Parameters.scala 121:31]
  wire [32:0] _T_127; // @[Parameters.scala 121:49]
  wire [32:0] _T_129; // @[Parameters.scala 121:52]
  wire  _T_130; // @[Parameters.scala 121:67]
  wire  _T_131; // @[Parameters.scala 168:56]
  wire [31:0] _T_133; // @[Parameters.scala 121:31]
  wire [32:0] _T_134; // @[Parameters.scala 121:49]
  wire [32:0] _T_136; // @[Parameters.scala 121:52]
  wire  _T_137; // @[Parameters.scala 121:67]
  wire [31:0] _T_138; // @[Parameters.scala 121:31]
  wire [32:0] _T_139; // @[Parameters.scala 121:49]
  wire [32:0] _T_141; // @[Parameters.scala 121:52]
  wire  _T_142; // @[Parameters.scala 121:67]
  wire [31:0] _T_143; // @[Parameters.scala 121:31]
  wire [32:0] _T_144; // @[Parameters.scala 121:49]
  wire [32:0] _T_146; // @[Parameters.scala 121:52]
  wire  _T_147; // @[Parameters.scala 121:67]
  wire [32:0] _T_151; // @[Parameters.scala 121:52]
  wire  _T_152; // @[Parameters.scala 121:67]
  wire [31:0] _T_153; // @[Parameters.scala 121:31]
  wire [32:0] _T_154; // @[Parameters.scala 121:49]
  wire [32:0] _T_156; // @[Parameters.scala 121:52]
  wire  _T_157; // @[Parameters.scala 121:67]
  wire [31:0] _T_158; // @[Parameters.scala 121:31]
  wire [32:0] _T_159; // @[Parameters.scala 121:49]
  wire [32:0] _T_161; // @[Parameters.scala 121:52]
  wire  _T_162; // @[Parameters.scala 121:67]
  wire  _T_163; // @[Parameters.scala 169:42]
  wire  _T_164; // @[Parameters.scala 169:42]
  wire  _T_165; // @[Parameters.scala 169:42]
  wire  _T_172; // @[Monitor.scala 49:14]
  wire  _T_184; // @[Parameters.scala 89:48]
  wire  _T_186; // @[Mux.scala 19:72]
  wire  _T_192; // @[Monitor.scala 50:14]
  wire  _T_195; // @[Monitor.scala 51:14]
  wire  _T_199; // @[Monitor.scala 52:14]
  wire  _T_202; // @[Monitor.scala 53:14]
  wire  _T_204; // @[Bundles.scala 109:27]
  wire  _T_206; // @[Monitor.scala 54:14]
  wire  _T_209; // @[Monitor.scala 55:28]
  wire  _T_211; // @[Monitor.scala 55:14]
  wire  _T_217; // @[Monitor.scala 59:25]
  wire  _T_304; // @[Monitor.scala 66:28]
  wire  _T_306; // @[Monitor.scala 66:14]
  wire  _T_317; // @[Monitor.scala 71:25]
  wire  _T_319; // @[Parameters.scala 90:42]
  wire  _T_327; // @[Parameters.scala 168:56]
  wire  _T_362; // @[Parameters.scala 169:42]
  wire  _T_363; // @[Parameters.scala 169:42]
  wire  _T_364; // @[Parameters.scala 169:42]
  wire  _T_365; // @[Parameters.scala 169:42]
  wire  _T_366; // @[Parameters.scala 169:42]
  wire  _T_367; // @[Parameters.scala 168:56]
  wire  _T_369; // @[Parameters.scala 170:30]
  wire  _T_371; // @[Monitor.scala 72:14]
  wire  _T_379; // @[Monitor.scala 75:28]
  wire  _T_381; // @[Monitor.scala 75:14]
  wire  _T_383; // @[Monitor.scala 76:27]
  wire  _T_385; // @[Monitor.scala 76:14]
  wire  _T_391; // @[Monitor.scala 80:25]
  wire  _T_428; // @[Parameters.scala 169:42]
  wire  _T_429; // @[Parameters.scala 168:56]
  wire  _T_431; // @[Parameters.scala 90:42]
  wire  _T_439; // @[Parameters.scala 168:56]
  wire  _T_448; // @[Parameters.scala 170:30]
  wire  _T_449; // @[Parameters.scala 170:30]
  wire  _T_452; // @[Monitor.scala 81:14]
  wire  _T_468; // @[Monitor.scala 88:25]
  wire [7:0] _T_542; // @[Monitor.scala 93:28]
  wire  _T_543; // @[Monitor.scala 93:37]
  wire  _T_545; // @[Monitor.scala 93:14]
  wire  _T_547; // @[Monitor.scala 96:25]
  wire  _T_549; // @[Parameters.scala 90:42]
  wire  _T_575; // @[Parameters.scala 168:56]
  wire  _T_598; // @[Monitor.scala 97:14]
  wire  _T_606; // @[Bundles.scala 139:33]
  wire  _T_608; // @[Monitor.scala 100:14]
  wire  _T_614; // @[Monitor.scala 104:25]
  wire  _T_673; // @[Bundles.scala 146:30]
  wire  _T_675; // @[Monitor.scala 108:14]
  wire  _T_681; // @[Monitor.scala 112:25]
  wire  _T_732; // @[Monitor.scala 113:14]
  wire  _T_748; // @[Bundles.scala 43:24]
  wire  _T_750; // @[Monitor.scala 268:12]
  wire  _T_762; // @[Parameters.scala 280:46]
  wire  _T_764; // @[Monitor.scala 275:25]
  wire  _T_766; // @[Monitor.scala 276:14]
  wire  _T_768; // @[Monitor.scala 277:27]
  wire  _T_770; // @[Monitor.scala 277:14]
  wire  _T_772; // @[Monitor.scala 278:28]
  wire  _T_774; // @[Monitor.scala 278:14]
  wire  _T_778; // @[Monitor.scala 279:14]
  wire  _T_782; // @[Monitor.scala 280:14]
  wire  _T_784; // @[Monitor.scala 283:25]
  wire  _T_795; // @[Bundles.scala 103:26]
  wire  _T_797; // @[Monitor.scala 287:14]
  wire  _T_799; // @[Monitor.scala 288:28]
  wire  _T_801; // @[Monitor.scala 288:14]
  wire  _T_812; // @[Monitor.scala 293:25]
  wire  _T_832; // @[Monitor.scala 299:30]
  wire  _T_834; // @[Monitor.scala 299:14]
  wire  _T_841; // @[Monitor.scala 303:25]
  wire  _T_858; // @[Monitor.scala 311:25]
  wire  _T_876; // @[Monitor.scala 319:25]
  wire  _T_893; // @[Bundles.scala 41:24]
  wire  _T_895; // @[Monitor.scala 122:12]
  wire [32:0] _T_900; // @[Parameters.scala 121:49]
  wire [31:0] _T_917; // @[Parameters.scala 121:31]
  wire [32:0] _T_918; // @[Parameters.scala 121:49]
  wire [32:0] _T_920; // @[Parameters.scala 121:52]
  wire  _T_921; // @[Parameters.scala 121:67]
  wire [31:0] _T_922; // @[Parameters.scala 121:31]
  wire [32:0] _T_923; // @[Parameters.scala 121:49]
  wire [32:0] _T_925; // @[Parameters.scala 121:52]
  wire  _T_926; // @[Parameters.scala 121:67]
  wire [31:0] _T_927; // @[Parameters.scala 121:31]
  wire [32:0] _T_928; // @[Parameters.scala 121:49]
  wire [32:0] _T_930; // @[Parameters.scala 121:52]
  wire  _T_931; // @[Parameters.scala 121:67]
  wire [32:0] _T_935; // @[Parameters.scala 121:52]
  wire  _T_936; // @[Parameters.scala 121:67]
  wire [31:0] _T_937; // @[Parameters.scala 121:31]
  wire [32:0] _T_938; // @[Parameters.scala 121:49]
  wire [32:0] _T_940; // @[Parameters.scala 121:52]
  wire  _T_941; // @[Parameters.scala 121:67]
  wire [31:0] _T_942; // @[Parameters.scala 121:31]
  wire [32:0] _T_943; // @[Parameters.scala 121:49]
  wire [32:0] _T_945; // @[Parameters.scala 121:52]
  wire  _T_946; // @[Parameters.scala 121:67]
  wire [31:0] _T_947; // @[Parameters.scala 121:31]
  wire [32:0] _T_948; // @[Parameters.scala 121:49]
  wire [32:0] _T_950; // @[Parameters.scala 121:52]
  wire  _T_951; // @[Parameters.scala 121:67]
  wire  _T_965; // @[Parameters.scala 155:64]
  wire  _T_966; // @[Parameters.scala 155:64]
  wire  _T_967; // @[Parameters.scala 155:64]
  wire  _T_968; // @[Parameters.scala 155:64]
  wire  _T_969; // @[Parameters.scala 155:64]
  wire  _T_970; // @[Parameters.scala 155:64]
  wire [26:0] _T_972; // @[package.scala 185:77]
  wire [31:0] _GEN_34; // @[Edges.scala 21:16]
  wire [31:0] _T_975; // @[Edges.scala 21:16]
  wire  _T_976; // @[Edges.scala 21:24]
  wire [3:0] _T_979; // @[OneHot.scala 52:12]
  wire [2:0] _T_981; // @[Misc.scala 206:81]
  wire  _T_982; // @[Misc.scala 210:21]
  wire  _T_987; // @[Misc.scala 219:38]
  wire  _T_988; // @[Misc.scala 219:29]
  wire  _T_990; // @[Misc.scala 219:38]
  wire  _T_991; // @[Misc.scala 219:29]
  wire  _T_995; // @[Misc.scala 218:27]
  wire  _T_996; // @[Misc.scala 219:38]
  wire  _T_997; // @[Misc.scala 219:29]
  wire  _T_998; // @[Misc.scala 218:27]
  wire  _T_999; // @[Misc.scala 219:38]
  wire  _T_1000; // @[Misc.scala 219:29]
  wire  _T_1001; // @[Misc.scala 218:27]
  wire  _T_1002; // @[Misc.scala 219:38]
  wire  _T_1003; // @[Misc.scala 219:29]
  wire  _T_1004; // @[Misc.scala 218:27]
  wire  _T_1005; // @[Misc.scala 219:38]
  wire  _T_1006; // @[Misc.scala 219:29]
  wire  _T_1010; // @[Misc.scala 218:27]
  wire  _T_1011; // @[Misc.scala 219:38]
  wire  _T_1012; // @[Misc.scala 219:29]
  wire  _T_1013; // @[Misc.scala 218:27]
  wire  _T_1014; // @[Misc.scala 219:38]
  wire  _T_1015; // @[Misc.scala 219:29]
  wire  _T_1016; // @[Misc.scala 218:27]
  wire  _T_1017; // @[Misc.scala 219:38]
  wire  _T_1018; // @[Misc.scala 219:29]
  wire  _T_1019; // @[Misc.scala 218:27]
  wire  _T_1020; // @[Misc.scala 219:38]
  wire  _T_1021; // @[Misc.scala 219:29]
  wire  _T_1022; // @[Misc.scala 218:27]
  wire  _T_1023; // @[Misc.scala 219:38]
  wire  _T_1024; // @[Misc.scala 219:29]
  wire  _T_1025; // @[Misc.scala 218:27]
  wire  _T_1026; // @[Misc.scala 219:38]
  wire  _T_1027; // @[Misc.scala 219:29]
  wire  _T_1028; // @[Misc.scala 218:27]
  wire  _T_1029; // @[Misc.scala 219:38]
  wire  _T_1030; // @[Misc.scala 219:29]
  wire  _T_1031; // @[Misc.scala 218:27]
  wire  _T_1032; // @[Misc.scala 219:38]
  wire  _T_1033; // @[Misc.scala 219:29]
  wire [7:0] _T_1040; // @[Cat.scala 30:58]
  wire  _T_1057; // @[Monitor.scala 130:117]
  wire  _T_1058; // @[Monitor.scala 132:25]
  wire  _T_1069; // @[Parameters.scala 89:48]
  wire  _T_1071; // @[Mux.scala 19:72]
  wire  _T_1077; // @[Monitor.scala 133:14]
  wire  _T_1080; // @[Monitor.scala 134:14]
  wire  _T_1083; // @[Monitor.scala 135:14]
  wire  _T_1086; // @[Monitor.scala 136:14]
  wire  _T_1088; // @[Bundles.scala 103:26]
  wire  _T_1090; // @[Monitor.scala 137:14]
  wire  _T_1092; // @[Monitor.scala 138:27]
  wire  _T_1094; // @[Monitor.scala 138:14]
  wire  _T_1098; // @[Monitor.scala 139:14]
  wire  _T_1100; // @[Monitor.scala 142:25]
  wire  _T_1113; // @[Monitor.scala 147:28]
  wire  _T_1115; // @[Monitor.scala 147:14]
  wire  _T_1125; // @[Monitor.scala 152:25]
  wire  _T_1146; // @[Monitor.scala 161:25]
  wire [7:0] _T_1164; // @[Monitor.scala 167:28]
  wire  _T_1165; // @[Monitor.scala 167:37]
  wire  _T_1167; // @[Monitor.scala 167:14]
  wire  _T_1169; // @[Monitor.scala 170:25]
  wire  _T_1190; // @[Monitor.scala 179:25]
  wire  _T_1211; // @[Monitor.scala 188:25]
  wire  _T_1246; // @[Parameters.scala 280:46]
  wire [26:0] _T_1248; // @[package.scala 185:77]
  wire [31:0] _GEN_35; // @[Edges.scala 21:16]
  wire [31:0] _T_1251; // @[Edges.scala 21:16]
  wire  _T_1252; // @[Edges.scala 21:24]
  wire [31:0] _T_1253; // @[Parameters.scala 121:31]
  wire [32:0] _T_1254; // @[Parameters.scala 121:49]
  wire [32:0] _T_1256; // @[Parameters.scala 121:52]
  wire  _T_1257; // @[Parameters.scala 121:67]
  wire [31:0] _T_1258; // @[Parameters.scala 121:31]
  wire [32:0] _T_1259; // @[Parameters.scala 121:49]
  wire [32:0] _T_1261; // @[Parameters.scala 121:52]
  wire  _T_1262; // @[Parameters.scala 121:67]
  wire [31:0] _T_1263; // @[Parameters.scala 121:31]
  wire [32:0] _T_1264; // @[Parameters.scala 121:49]
  wire [32:0] _T_1266; // @[Parameters.scala 121:52]
  wire  _T_1267; // @[Parameters.scala 121:67]
  wire [32:0] _T_1269; // @[Parameters.scala 121:49]
  wire [32:0] _T_1271; // @[Parameters.scala 121:52]
  wire  _T_1272; // @[Parameters.scala 121:67]
  wire [31:0] _T_1273; // @[Parameters.scala 121:31]
  wire [32:0] _T_1274; // @[Parameters.scala 121:49]
  wire [32:0] _T_1276; // @[Parameters.scala 121:52]
  wire  _T_1277; // @[Parameters.scala 121:67]
  wire [31:0] _T_1278; // @[Parameters.scala 121:31]
  wire [32:0] _T_1279; // @[Parameters.scala 121:49]
  wire [32:0] _T_1281; // @[Parameters.scala 121:52]
  wire  _T_1282; // @[Parameters.scala 121:67]
  wire [31:0] _T_1283; // @[Parameters.scala 121:31]
  wire [32:0] _T_1284; // @[Parameters.scala 121:49]
  wire [32:0] _T_1286; // @[Parameters.scala 121:52]
  wire  _T_1287; // @[Parameters.scala 121:67]
  wire  _T_1301; // @[Parameters.scala 155:64]
  wire  _T_1302; // @[Parameters.scala 155:64]
  wire  _T_1303; // @[Parameters.scala 155:64]
  wire  _T_1304; // @[Parameters.scala 155:64]
  wire  _T_1305; // @[Parameters.scala 155:64]
  wire  _T_1306; // @[Parameters.scala 155:64]
  wire  _T_1327; // @[Monitor.scala 207:25]
  wire  _T_1329; // @[Monitor.scala 208:14]
  wire  _T_1332; // @[Monitor.scala 209:14]
  wire  _T_1334; // @[Monitor.scala 210:27]
  wire  _T_1336; // @[Monitor.scala 210:14]
  wire  _T_1339; // @[Monitor.scala 211:14]
  wire  _T_1341; // @[Bundles.scala 121:29]
  wire  _T_1343; // @[Monitor.scala 212:14]
  wire  _T_1349; // @[Monitor.scala 216:25]
  wire  _T_1367; // @[Monitor.scala 224:25]
  wire  _T_1369; // @[Parameters.scala 90:42]
  wire  _T_1377; // @[Parameters.scala 168:56]
  wire  _T_1418; // @[Monitor.scala 225:14]
  wire  _T_1430; // @[Parameters.scala 89:48]
  wire  _T_1432; // @[Mux.scala 19:72]
  wire  _T_1438; // @[Monitor.scala 226:14]
  wire  _T_1450; // @[Bundles.scala 115:29]
  wire  _T_1452; // @[Monitor.scala 230:14]
  wire  _T_1458; // @[Monitor.scala 234:25]
  wire  _T_1545; // @[Monitor.scala 243:25]
  wire  _T_1555; // @[Monitor.scala 247:28]
  wire  _T_1557; // @[Monitor.scala 247:14]
  wire  _T_1563; // @[Monitor.scala 251:25]
  wire  _T_1577; // @[Monitor.scala 258:25]
  wire  _T_1599; // @[Bundles.scala 277:22]
  wire [8:0] _T_1604; // @[Edges.scala 220:59]
  reg [8:0] _T_1609; // @[Edges.scala 229:27]
  reg [31:0] _RAND_0;
  wire [8:0] _T_1612; // @[Edges.scala 230:28]
  wire  _T_1613; // @[Edges.scala 231:25]
  reg [2:0] _T_1622; // @[Monitor.scala 349:22]
  reg [31:0] _RAND_1;
  reg [2:0] _T_1624; // @[Monitor.scala 350:22]
  reg [31:0] _RAND_2;
  reg [3:0] _T_1626; // @[Monitor.scala 351:22]
  reg [31:0] _RAND_3;
  reg  _T_1628; // @[Monitor.scala 352:22]
  reg [31:0] _RAND_4;
  reg [31:0] _T_1630; // @[Monitor.scala 353:22]
  reg [31:0] _RAND_5;
  wire  _T_1632; // @[Monitor.scala 354:19]
  wire  _T_1633; // @[Monitor.scala 355:29]
  wire  _T_1635; // @[Monitor.scala 355:14]
  wire  _T_1637; // @[Monitor.scala 356:29]
  wire  _T_1639; // @[Monitor.scala 356:14]
  wire  _T_1641; // @[Monitor.scala 357:29]
  wire  _T_1643; // @[Monitor.scala 357:14]
  wire  _T_1645; // @[Monitor.scala 358:29]
  wire  _T_1647; // @[Monitor.scala 358:14]
  wire  _T_1649; // @[Monitor.scala 359:29]
  wire  _T_1651; // @[Monitor.scala 359:14]
  wire  _T_1654; // @[Monitor.scala 361:20]
  wire  _T_1655; // @[Bundles.scala 277:22]
  wire [26:0] _T_1657; // @[package.scala 185:77]
  wire [8:0] _T_1660; // @[Edges.scala 220:59]
  reg [8:0] _T_1664; // @[Edges.scala 229:27]
  reg [31:0] _RAND_6;
  wire [8:0] _T_1667; // @[Edges.scala 230:28]
  wire  _T_1668; // @[Edges.scala 231:25]
  reg [2:0] _T_1677; // @[Monitor.scala 418:22]
  reg [31:0] _RAND_7;
  reg [1:0] _T_1679; // @[Monitor.scala 419:22]
  reg [31:0] _RAND_8;
  reg [3:0] _T_1681; // @[Monitor.scala 420:22]
  reg [31:0] _RAND_9;
  reg  _T_1683; // @[Monitor.scala 421:22]
  reg [31:0] _RAND_10;
  reg [1:0] _T_1685; // @[Monitor.scala 422:22]
  reg [31:0] _RAND_11;
  reg  _T_1687; // @[Monitor.scala 423:22]
  reg [31:0] _RAND_12;
  wire  _T_1689; // @[Monitor.scala 424:19]
  wire  _T_1690; // @[Monitor.scala 425:29]
  wire  _T_1692; // @[Monitor.scala 425:14]
  wire  _T_1694; // @[Monitor.scala 426:29]
  wire  _T_1696; // @[Monitor.scala 426:14]
  wire  _T_1698; // @[Monitor.scala 427:29]
  wire  _T_1700; // @[Monitor.scala 427:14]
  wire  _T_1702; // @[Monitor.scala 428:29]
  wire  _T_1704; // @[Monitor.scala 428:14]
  wire  _T_1706; // @[Monitor.scala 429:29]
  wire  _T_1708; // @[Monitor.scala 429:14]
  wire  _T_1710; // @[Monitor.scala 430:29]
  wire  _T_1712; // @[Monitor.scala 430:14]
  wire  _T_1715; // @[Monitor.scala 432:20]
  wire  _T_1716; // @[Bundles.scala 277:22]
  reg [8:0] _T_1726; // @[Edges.scala 229:27]
  reg [31:0] _RAND_13;
  wire [8:0] _T_1729; // @[Edges.scala 230:28]
  wire  _T_1730; // @[Edges.scala 231:25]
  reg [2:0] _T_1739; // @[Monitor.scala 372:22]
  reg [31:0] _RAND_14;
  reg [1:0] _T_1741; // @[Monitor.scala 373:22]
  reg [31:0] _RAND_15;
  reg [3:0] _T_1743; // @[Monitor.scala 374:22]
  reg [31:0] _RAND_16;
  reg  _T_1745; // @[Monitor.scala 375:22]
  reg [31:0] _RAND_17;
  reg [31:0] _T_1747; // @[Monitor.scala 376:22]
  reg [31:0] _RAND_18;
  wire  _T_1749; // @[Monitor.scala 377:19]
  wire  _T_1750; // @[Monitor.scala 378:29]
  wire  _T_1752; // @[Monitor.scala 378:14]
  wire  _T_1754; // @[Monitor.scala 379:29]
  wire  _T_1756; // @[Monitor.scala 379:14]
  wire  _T_1758; // @[Monitor.scala 380:29]
  wire  _T_1760; // @[Monitor.scala 380:14]
  wire  _T_1762; // @[Monitor.scala 381:29]
  wire  _T_1764; // @[Monitor.scala 381:14]
  wire  _T_1766; // @[Monitor.scala 382:29]
  wire  _T_1768; // @[Monitor.scala 382:14]
  wire  _T_1771; // @[Monitor.scala 384:20]
  wire  _T_1772; // @[Bundles.scala 277:22]
  wire [8:0] _T_1777; // @[Edges.scala 220:59]
  reg [8:0] _T_1781; // @[Edges.scala 229:27]
  reg [31:0] _RAND_19;
  wire [8:0] _T_1784; // @[Edges.scala 230:28]
  wire  _T_1785; // @[Edges.scala 231:25]
  reg [2:0] _T_1794; // @[Monitor.scala 395:22]
  reg [31:0] _RAND_20;
  reg [2:0] _T_1796; // @[Monitor.scala 396:22]
  reg [31:0] _RAND_21;
  reg [3:0] _T_1798; // @[Monitor.scala 397:22]
  reg [31:0] _RAND_22;
  reg  _T_1800; // @[Monitor.scala 398:22]
  reg [31:0] _RAND_23;
  reg [31:0] _T_1802; // @[Monitor.scala 399:22]
  reg [31:0] _RAND_24;
  wire  _T_1804; // @[Monitor.scala 400:19]
  wire  _T_1805; // @[Monitor.scala 401:29]
  wire  _T_1807; // @[Monitor.scala 401:14]
  wire  _T_1809; // @[Monitor.scala 402:29]
  wire  _T_1811; // @[Monitor.scala 402:14]
  wire  _T_1813; // @[Monitor.scala 403:29]
  wire  _T_1815; // @[Monitor.scala 403:14]
  wire  _T_1817; // @[Monitor.scala 404:29]
  wire  _T_1819; // @[Monitor.scala 404:14]
  wire  _T_1821; // @[Monitor.scala 405:29]
  wire  _T_1823; // @[Monitor.scala 405:14]
  wire  _T_1826; // @[Monitor.scala 407:20]
  reg [1:0] _T_1828; // @[Monitor.scala 452:27]
  reg [31:0] _RAND_25;
  reg [8:0] _T_1839; // @[Edges.scala 229:27]
  reg [31:0] _RAND_26;
  wire [8:0] _T_1842; // @[Edges.scala 230:28]
  wire  _T_1843; // @[Edges.scala 231:25]
  reg [8:0] _T_1860; // @[Edges.scala 229:27]
  reg [31:0] _RAND_27;
  wire [8:0] _T_1863; // @[Edges.scala 230:28]
  wire  _T_1864; // @[Edges.scala 231:25]
  wire  _T_1875; // @[Monitor.scala 458:27]
  wire [1:0] _T_1877; // @[OneHot.scala 45:35]
  wire [1:0] _T_1878; // @[Monitor.scala 460:23]
  wire  _T_1882; // @[Monitor.scala 460:13]
  wire [1:0] _GEN_27; // @[Monitor.scala 458:72]
  wire  _T_1888; // @[Monitor.scala 465:27]
  wire  _T_1891; // @[Monitor.scala 465:72]
  wire [1:0] _T_1892; // @[OneHot.scala 45:35]
  wire [1:0] _T_1893; // @[Monitor.scala 467:21]
  wire [1:0] _T_1894; // @[Monitor.scala 467:32]
  wire  _T_1897; // @[Monitor.scala 467:13]
  wire [1:0] _GEN_28; // @[Monitor.scala 465:91]
  wire  _T_1899; // @[Monitor.scala 471:20]
  wire  _T_1900; // @[Monitor.scala 471:40]
  wire  _T_1902; // @[Monitor.scala 471:30]
  wire  _T_1904; // @[Monitor.scala 471:13]
  wire [1:0] _T_1906; // @[Monitor.scala 474:27]
  wire [1:0] _T_1908; // @[Monitor.scala 474:36]
  reg [3:0] _T_1926; // @[Monitor.scala 486:27]
  reg [31:0] _RAND_28;
  reg [8:0] _T_1936; // @[Edges.scala 229:27]
  reg [31:0] _RAND_29;
  wire [8:0] _T_1939; // @[Edges.scala 230:28]
  wire  _T_1940; // @[Edges.scala 231:25]
  wire  _T_1951; // @[Monitor.scala 492:27]
  wire  _T_1955; // @[Edges.scala 71:40]
  wire  _T_1956; // @[Monitor.scala 492:38]
  wire [3:0] _T_1957; // @[OneHot.scala 45:35]
  wire [3:0] _T_1958; // @[Monitor.scala 494:23]
  wire  _T_1962; // @[Monitor.scala 494:13]
  wire [3:0] _GEN_31; // @[Monitor.scala 492:72]
  wire  _T_1966; // @[Bundles.scala 277:22]
  wire [3:0] _T_1969; // @[OneHot.scala 45:35]
  wire [3:0] _T_1970; // @[Monitor.scala 500:21]
  wire [3:0] _T_1971; // @[Monitor.scala 500:32]
  wire  _T_1974; // @[Monitor.scala 500:13]
  wire [3:0] _GEN_32; // @[Monitor.scala 498:73]
  wire [3:0] _T_1976; // @[Monitor.scala 505:27]
  wire [3:0] _T_1978; // @[Monitor.scala 505:36]
  wire  _GEN_36; // @[Monitor.scala 49:14]
  wire  _GEN_50; // @[Monitor.scala 60:14]
  wire  _GEN_66; // @[Monitor.scala 72:14]
  wire  _GEN_76; // @[Monitor.scala 81:14]
  wire  _GEN_86; // @[Monitor.scala 89:14]
  wire  _GEN_96; // @[Monitor.scala 97:14]
  wire  _GEN_106; // @[Monitor.scala 105:14]
  wire  _GEN_116; // @[Monitor.scala 113:14]
  wire  _GEN_124; // @[Monitor.scala 276:14]
  wire  _GEN_134; // @[Monitor.scala 284:14]
  wire  _GEN_144; // @[Monitor.scala 294:14]
  wire  _GEN_154; // @[Monitor.scala 304:14]
  wire  _GEN_160; // @[Monitor.scala 312:14]
  wire  _GEN_166; // @[Monitor.scala 320:14]
  wire  _GEN_172; // @[Monitor.scala 133:14]
  wire  _GEN_186; // @[Monitor.scala 143:14]
  wire  _GEN_200; // @[Monitor.scala 153:14]
  wire  _GEN_212; // @[Monitor.scala 162:14]
  wire  _GEN_224; // @[Monitor.scala 171:14]
  wire  _GEN_234; // @[Monitor.scala 180:14]
  wire  _GEN_244; // @[Monitor.scala 189:14]
  wire  _GEN_256; // @[Monitor.scala 208:14]
  wire  _GEN_266; // @[Monitor.scala 217:14]
  wire  _GEN_276; // @[Monitor.scala 225:14]
  wire  _GEN_288; // @[Monitor.scala 235:14]
  wire  _GEN_300; // @[Monitor.scala 244:14]
  wire  _GEN_308; // @[Monitor.scala 252:14]
  wire  _GEN_316; // @[Monitor.scala 259:14]
  wire [29:0] TLMonitor_64_covSum;
  wire  stopEn0;
  wire  stopEn1;
  wire  stopEn2;
  wire  stopEn3;
  wire  stopEn4;
  wire  stopEn5;
  wire  stopEn6;
  wire  stopEn7;
  wire  stopEn8;
  wire  stopEn9;
  wire  stopEn10;
  wire  stopEn11;
  wire  stopEn12;
  wire  stopEn13;
  wire  stopEn14;
  wire  stopEn15;
  wire  stopEn16;
  wire  stopEn17;
  wire  stopEn18;
  wire  stopEn19;
  wire  stopEn20;
  wire  stopEn21;
  wire  stopEn22;
  wire  stopEn23;
  wire  stopEn24;
  wire  stopEn25;
  wire  stopEn26;
  wire  stopEn27;
  wire  stopEn28;
  wire  stopEn29;
  wire  stopEn30;
  wire  stopEn31;
  wire  stopEn32;
  wire  stopEn33;
  wire  stopEn34;
  wire  stopEn35;
  wire  stopEn36;
  wire  stopEn37;
  wire  stopEn38;
  wire  stopEn39;
  wire  stopEn40;
  wire  stopEn41;
  wire  stopEn42;
  wire  stopEn43;
  wire  stopEn44;
  wire  stopEn45;
  wire  stopEn46;
  wire  stopEn47;
  wire  stopEn48;
  wire  stopEn49;
  wire  stopEn50;
  wire  stopEn51;
  wire  stopEn52;
  wire  stopEn53;
  wire  stopEn54;
  wire  stopEn55;
  wire  stopEn56;
  wire  stopEn57;
  wire  stopEn58;
  wire  stopEn59;
  wire  stopEn60;
  wire  stopEn61;
  wire  stopEn62;
  wire  stopEn63;
  wire  stopEn64;
  wire  stopEn65;
  wire  stopEn66;
  wire  stopEn67;
  wire  stopEn68;
  wire  stopEn69;
  wire  stopEn70;
  wire  stopEn71;
  wire  stopEn72;
  wire  stopEn73;
  wire  stopEn74;
  wire  stopEn75;
  wire  stopEn76;
  wire  stopEn77;
  wire  stopEn78;
  wire  stopEn79;
  wire  stopEn80;
  wire  stopEn81;
  wire  stopEn82;
  wire  stopEn83;
  wire  stopEn84;
  wire  stopEn85;
  wire  stopEn86;
  wire  stopEn87;
  wire  stopEn88;
  wire  stopEn89;
  wire  stopEn90;
  wire  stopEn91;
  wire  stopEn92;
  wire  stopEn93;
  wire  stopEn94;
  wire  stopEn95;
  wire  stopEn96;
  wire  stopEn97;
  wire  stopEn98;
  wire  stopEn99;
  wire  stopEn100;
  wire  stopEn101;
  wire  stopEn102;
  wire  stopEn103;
  wire  stopEn104;
  wire  stopEn105;
  wire  stopEn106;
  wire  stopEn107;
  wire  stopEn108;
  wire  stopEn109;
  wire  stopEn110;
  wire  stopEn111;
  wire  stopEn112;
  wire  stopEn113;
  wire  stopEn114;
  wire  stopEn115;
  wire  stopEn116;
  wire  stopEn117;
  wire  stopEn118;
  wire  stopEn119;
  wire  stopEn120;
  wire  stopEn121;
  wire  stopEn122;
  wire  stopEn123;
  wire  stopEn124;
  wire  stopEn125;
  wire  stopEn126;
  wire  stopEn127;
  wire  stopEn128;
  wire  stopEn129;
  wire  stopEn130;
  wire  stopEn131;
  wire  stopEn132;
  wire  stopEn133;
  wire  stopEn134;
  wire  stopEn135;
  wire  stopEn136;
  wire  stopEn137;
  wire  stopEn138;
  wire  stopEn139;
  wire  stopEn140;
  wire  stopEn141;
  wire  stopEn142;
  wire  stopEn143;
  wire  stopEn144;
  wire  stopEn145;
  wire  stopEn146;
  wire  stopEn147;
  wire  stopEn148;
  wire  stopEn149;
  wire  stopEn150;
  wire  stopEn151;
  wire  stopEn152;
  wire  stopEn153;
  wire  stopEn154;
  wire  stopEn155;
  wire  stopEn156;
  wire  stopEn157;
  wire  stopEn158;
  wire  stopEn159;
  wire  stopEn160;
  wire  stopEn161;
  wire  stopEn162;
  wire  stopEn163;
  wire  stopEn164;
  wire  stopEn165;
  wire  stopEn166;
  wire  stopEn167;
  wire  stopEn168;
  wire  stopEn169;
  wire  stopEn170;
  wire  stopEn171;
  wire  TLMonitor_64_or63;
  wire  TLMonitor_64_or130;
  wire  TLMonitor_64_or64;
  wire  TLMonitor_64_or31;
  wire  TLMonitor_64_or65;
  wire  TLMonitor_64_or134;
  wire  TLMonitor_64_or66;
  wire  TLMonitor_64_or32;
  wire  TLMonitor_64_or15;
  wire  TLMonitor_64_or67;
  wire  TLMonitor_64_or138;
  wire  TLMonitor_64_or68;
  wire  TLMonitor_64_or33;
  wire  TLMonitor_64_or140;
  wire  TLMonitor_64_or69;
  wire  TLMonitor_64_or142;
  wire  TLMonitor_64_or70;
  wire  TLMonitor_64_or34;
  wire  TLMonitor_64_or16;
  wire  TLMonitor_64_or7;
  wire  TLMonitor_64_or71;
  wire  TLMonitor_64_or146;
  wire  TLMonitor_64_or72;
  wire  TLMonitor_64_or35;
  wire  TLMonitor_64_or148;
  wire  TLMonitor_64_or73;
  wire  TLMonitor_64_or150;
  wire  TLMonitor_64_or74;
  wire  TLMonitor_64_or36;
  wire  TLMonitor_64_or17;
  wire  TLMonitor_64_or75;
  wire  TLMonitor_64_or154;
  wire  TLMonitor_64_or76;
  wire  TLMonitor_64_or37;
  wire  TLMonitor_64_or156;
  wire  TLMonitor_64_or77;
  wire  TLMonitor_64_or158;
  wire  TLMonitor_64_or78;
  wire  TLMonitor_64_or38;
  wire  TLMonitor_64_or18;
  wire  TLMonitor_64_or8;
  wire  TLMonitor_64_or3;
  wire  TLMonitor_64_or79;
  wire  TLMonitor_64_or162;
  wire  TLMonitor_64_or80;
  wire  TLMonitor_64_or39;
  wire  TLMonitor_64_or81;
  wire  TLMonitor_64_or166;
  wire  TLMonitor_64_or82;
  wire  TLMonitor_64_or40;
  wire  TLMonitor_64_or19;
  wire  TLMonitor_64_or83;
  wire  TLMonitor_64_or170;
  wire  TLMonitor_64_or84;
  wire  TLMonitor_64_or41;
  wire  TLMonitor_64_or172;
  wire  TLMonitor_64_or85;
  wire  TLMonitor_64_or174;
  wire  TLMonitor_64_or86;
  wire  TLMonitor_64_or42;
  wire  TLMonitor_64_or20;
  wire  TLMonitor_64_or9;
  wire  TLMonitor_64_or87;
  wire  TLMonitor_64_or178;
  wire  TLMonitor_64_or88;
  wire  TLMonitor_64_or43;
  wire  TLMonitor_64_or180;
  wire  TLMonitor_64_or89;
  wire  TLMonitor_64_or182;
  wire  TLMonitor_64_or90;
  wire  TLMonitor_64_or44;
  wire  TLMonitor_64_or21;
  wire  TLMonitor_64_or91;
  wire  TLMonitor_64_or186;
  wire  TLMonitor_64_or92;
  wire  TLMonitor_64_or45;
  wire  TLMonitor_64_or188;
  wire  TLMonitor_64_or93;
  wire  TLMonitor_64_or190;
  wire  TLMonitor_64_or94;
  wire  TLMonitor_64_or46;
  wire  TLMonitor_64_or22;
  wire  TLMonitor_64_or10;
  wire  TLMonitor_64_or4;
  wire  TLMonitor_64_or1;
  wire  TLMonitor_64_or95;
  wire  TLMonitor_64_or194;
  wire  TLMonitor_64_or96;
  wire  TLMonitor_64_or47;
  wire  TLMonitor_64_or97;
  wire  TLMonitor_64_or198;
  wire  TLMonitor_64_or98;
  wire  TLMonitor_64_or48;
  wire  TLMonitor_64_or23;
  wire  TLMonitor_64_or99;
  wire  TLMonitor_64_or202;
  wire  TLMonitor_64_or100;
  wire  TLMonitor_64_or49;
  wire  TLMonitor_64_or204;
  wire  TLMonitor_64_or101;
  wire  TLMonitor_64_or206;
  wire  TLMonitor_64_or102;
  wire  TLMonitor_64_or50;
  wire  TLMonitor_64_or24;
  wire  TLMonitor_64_or11;
  wire  TLMonitor_64_or103;
  wire  TLMonitor_64_or210;
  wire  TLMonitor_64_or104;
  wire  TLMonitor_64_or51;
  wire  TLMonitor_64_or212;
  wire  TLMonitor_64_or105;
  wire  TLMonitor_64_or214;
  wire  TLMonitor_64_or106;
  wire  TLMonitor_64_or52;
  wire  TLMonitor_64_or25;
  wire  TLMonitor_64_or107;
  wire  TLMonitor_64_or218;
  wire  TLMonitor_64_or108;
  wire  TLMonitor_64_or53;
  wire  TLMonitor_64_or220;
  wire  TLMonitor_64_or109;
  wire  TLMonitor_64_or222;
  wire  TLMonitor_64_or110;
  wire  TLMonitor_64_or54;
  wire  TLMonitor_64_or26;
  wire  TLMonitor_64_or12;
  wire  TLMonitor_64_or5;
  wire  TLMonitor_64_or111;
  wire  TLMonitor_64_or226;
  wire  TLMonitor_64_or112;
  wire  TLMonitor_64_or55;
  wire  TLMonitor_64_or113;
  wire  TLMonitor_64_or230;
  wire  TLMonitor_64_or114;
  wire  TLMonitor_64_or56;
  wire  TLMonitor_64_or27;
  wire  TLMonitor_64_or115;
  wire  TLMonitor_64_or234;
  wire  TLMonitor_64_or116;
  wire  TLMonitor_64_or57;
  wire  TLMonitor_64_or236;
  wire  TLMonitor_64_or117;
  wire  TLMonitor_64_or238;
  wire  TLMonitor_64_or118;
  wire  TLMonitor_64_or58;
  wire  TLMonitor_64_or28;
  wire  TLMonitor_64_or13;
  wire  TLMonitor_64_or119;
  wire  TLMonitor_64_or242;
  wire  TLMonitor_64_or120;
  wire  TLMonitor_64_or59;
  wire  TLMonitor_64_or244;
  wire  TLMonitor_64_or121;
  wire  TLMonitor_64_or246;
  wire  TLMonitor_64_or122;
  wire  TLMonitor_64_or60;
  wire  TLMonitor_64_or29;
  wire  TLMonitor_64_or123;
  wire  TLMonitor_64_or250;
  wire  TLMonitor_64_or124;
  wire  TLMonitor_64_or61;
  wire  TLMonitor_64_or252;
  wire  TLMonitor_64_or125;
  wire  TLMonitor_64_or254;
  wire  TLMonitor_64_or126;
  wire  TLMonitor_64_or62;
  wire  TLMonitor_64_or30;
  wire  TLMonitor_64_or14;
  wire  TLMonitor_64_or6;
  wire  TLMonitor_64_or2;
  wire  TLMonitor_64_or0;
  reg  TLMonitor_64_metaAssert;
  reg [31:0] _RAND_30;
  assign _T_30 = ~io_in_a_bits_source | io_in_a_bits_source; // @[Parameters.scala 280:46]
  assign _T_32 = 27'hfff << io_in_a_bits_size; // @[package.scala 185:77]
  assign _GEN_33 = {{20'd0}, ~_T_32[11:0]}; // @[Edges.scala 21:16]
  assign _T_35 = io_in_a_bits_address & _GEN_33; // @[Edges.scala 21:16]
  assign _T_36 = _T_35 == 32'h0; // @[Edges.scala 21:24]
  assign _T_39 = 4'h1 << io_in_a_bits_size[1:0]; // @[OneHot.scala 52:12]
  assign _T_41 = _T_39[2:0] | 3'h1; // @[Misc.scala 206:81]
  assign _T_42 = io_in_a_bits_size >= 4'h3; // @[Misc.scala 210:21]
  assign _T_47 = _T_41[2] & ~io_in_a_bits_address[2]; // @[Misc.scala 219:38]
  assign _T_48 = _T_42 | _T_47; // @[Misc.scala 219:29]
  assign _T_50 = _T_41[2] & io_in_a_bits_address[2]; // @[Misc.scala 219:38]
  assign _T_51 = _T_42 | _T_50; // @[Misc.scala 219:29]
  assign _T_55 = ~io_in_a_bits_address[2] & ~io_in_a_bits_address[1]; // @[Misc.scala 218:27]
  assign _T_56 = _T_41[1] & _T_55; // @[Misc.scala 219:38]
  assign _T_57 = _T_48 | _T_56; // @[Misc.scala 219:29]
  assign _T_58 = ~io_in_a_bits_address[2] & io_in_a_bits_address[1]; // @[Misc.scala 218:27]
  assign _T_59 = _T_41[1] & _T_58; // @[Misc.scala 219:38]
  assign _T_60 = _T_48 | _T_59; // @[Misc.scala 219:29]
  assign _T_61 = io_in_a_bits_address[2] & ~io_in_a_bits_address[1]; // @[Misc.scala 218:27]
  assign _T_62 = _T_41[1] & _T_61; // @[Misc.scala 219:38]
  assign _T_63 = _T_51 | _T_62; // @[Misc.scala 219:29]
  assign _T_64 = io_in_a_bits_address[2] & io_in_a_bits_address[1]; // @[Misc.scala 218:27]
  assign _T_65 = _T_41[1] & _T_64; // @[Misc.scala 219:38]
  assign _T_66 = _T_51 | _T_65; // @[Misc.scala 219:29]
  assign _T_70 = _T_55 & ~io_in_a_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_71 = _T_41[0] & _T_70; // @[Misc.scala 219:38]
  assign _T_72 = _T_57 | _T_71; // @[Misc.scala 219:29]
  assign _T_73 = _T_55 & io_in_a_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_74 = _T_41[0] & _T_73; // @[Misc.scala 219:38]
  assign _T_75 = _T_57 | _T_74; // @[Misc.scala 219:29]
  assign _T_76 = _T_58 & ~io_in_a_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_77 = _T_41[0] & _T_76; // @[Misc.scala 219:38]
  assign _T_78 = _T_60 | _T_77; // @[Misc.scala 219:29]
  assign _T_79 = _T_58 & io_in_a_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_80 = _T_41[0] & _T_79; // @[Misc.scala 219:38]
  assign _T_81 = _T_60 | _T_80; // @[Misc.scala 219:29]
  assign _T_82 = _T_61 & ~io_in_a_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_83 = _T_41[0] & _T_82; // @[Misc.scala 219:38]
  assign _T_84 = _T_63 | _T_83; // @[Misc.scala 219:29]
  assign _T_85 = _T_61 & io_in_a_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_86 = _T_41[0] & _T_85; // @[Misc.scala 219:38]
  assign _T_87 = _T_63 | _T_86; // @[Misc.scala 219:29]
  assign _T_88 = _T_64 & ~io_in_a_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_89 = _T_41[0] & _T_88; // @[Misc.scala 219:38]
  assign _T_90 = _T_66 | _T_89; // @[Misc.scala 219:29]
  assign _T_91 = _T_64 & io_in_a_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_92 = _T_41[0] & _T_91; // @[Misc.scala 219:38]
  assign _T_93 = _T_66 | _T_92; // @[Misc.scala 219:29]
  assign _T_100 = {_T_93,_T_90,_T_87,_T_84,_T_81,_T_78,_T_75,_T_72}; // @[Cat.scala 30:58]
  assign _T_104 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 121:49]
  assign _T_121 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 48:25]
  assign _T_123 = io_in_a_bits_size <= 4'h6; // @[Parameters.scala 90:42]
  assign _T_126 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 121:31]
  assign _T_127 = {1'b0,$signed(_T_126)}; // @[Parameters.scala 121:49]
  assign _T_129 = $signed(_T_127) & -33'sh10000000; // @[Parameters.scala 121:52]
  assign _T_130 = $signed(_T_129) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_131 = _T_123 & _T_130; // @[Parameters.scala 168:56]
  assign _T_133 = io_in_a_bits_address ^ 32'h3000; // @[Parameters.scala 121:31]
  assign _T_134 = {1'b0,$signed(_T_133)}; // @[Parameters.scala 121:49]
  assign _T_136 = $signed(_T_134) & -33'sh1000; // @[Parameters.scala 121:52]
  assign _T_137 = $signed(_T_136) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_138 = io_in_a_bits_address ^ 32'hc000000; // @[Parameters.scala 121:31]
  assign _T_139 = {1'b0,$signed(_T_138)}; // @[Parameters.scala 121:49]
  assign _T_141 = $signed(_T_139) & -33'sh4000000; // @[Parameters.scala 121:52]
  assign _T_142 = $signed(_T_141) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_143 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 121:31]
  assign _T_144 = {1'b0,$signed(_T_143)}; // @[Parameters.scala 121:49]
  assign _T_146 = $signed(_T_144) & -33'sh10000; // @[Parameters.scala 121:52]
  assign _T_147 = $signed(_T_146) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_151 = $signed(_T_104) & -33'sh1000; // @[Parameters.scala 121:52]
  assign _T_152 = $signed(_T_151) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_153 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 121:31]
  assign _T_154 = {1'b0,$signed(_T_153)}; // @[Parameters.scala 121:49]
  assign _T_156 = $signed(_T_154) & -33'sh10000; // @[Parameters.scala 121:52]
  assign _T_157 = $signed(_T_156) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_158 = io_in_a_bits_address ^ 32'h60000000; // @[Parameters.scala 121:31]
  assign _T_159 = {1'b0,$signed(_T_158)}; // @[Parameters.scala 121:49]
  assign _T_161 = $signed(_T_159) & -33'sh20000000; // @[Parameters.scala 121:52]
  assign _T_162 = $signed(_T_161) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_163 = _T_137 | _T_142; // @[Parameters.scala 169:42]
  assign _T_164 = _T_163 | _T_147; // @[Parameters.scala 169:42]
  assign _T_165 = _T_164 | _T_152; // @[Parameters.scala 169:42]
  assign _T_172 = _T_131 | reset; // @[Monitor.scala 49:14]
  assign _T_184 = 4'h6 == io_in_a_bits_size; // @[Parameters.scala 89:48]
  assign _T_186 = ~io_in_a_bits_source & _T_184; // @[Mux.scala 19:72]
  assign _T_192 = _T_186 | reset; // @[Monitor.scala 50:14]
  assign _T_195 = _T_30 | reset; // @[Monitor.scala 51:14]
  assign _T_199 = _T_42 | reset; // @[Monitor.scala 52:14]
  assign _T_202 = _T_36 | reset; // @[Monitor.scala 53:14]
  assign _T_204 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 109:27]
  assign _T_206 = _T_204 | reset; // @[Monitor.scala 54:14]
  assign _T_209 = ~io_in_a_bits_mask == 8'h0; // @[Monitor.scala 55:28]
  assign _T_211 = _T_209 | reset; // @[Monitor.scala 55:14]
  assign _T_217 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 59:25]
  assign _T_304 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 66:28]
  assign _T_306 = _T_304 | reset; // @[Monitor.scala 66:14]
  assign _T_317 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 71:25]
  assign _T_319 = io_in_a_bits_size <= 4'hc; // @[Parameters.scala 90:42]
  assign _T_327 = _T_319 & _T_137; // @[Parameters.scala 168:56]
  assign _T_362 = _T_142 | _T_147; // @[Parameters.scala 169:42]
  assign _T_363 = _T_362 | _T_152; // @[Parameters.scala 169:42]
  assign _T_364 = _T_363 | _T_157; // @[Parameters.scala 169:42]
  assign _T_365 = _T_364 | _T_130; // @[Parameters.scala 169:42]
  assign _T_366 = _T_365 | _T_162; // @[Parameters.scala 169:42]
  assign _T_367 = _T_123 & _T_366; // @[Parameters.scala 168:56]
  assign _T_369 = _T_327 | _T_367; // @[Parameters.scala 170:30]
  assign _T_371 = _T_369 | reset; // @[Monitor.scala 72:14]
  assign _T_379 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 75:28]
  assign _T_381 = _T_379 | reset; // @[Monitor.scala 75:14]
  assign _T_383 = io_in_a_bits_mask == _T_100; // @[Monitor.scala 76:27]
  assign _T_385 = _T_383 | reset; // @[Monitor.scala 76:14]
  assign _T_391 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 80:25]
  assign _T_428 = _T_363 | _T_130; // @[Parameters.scala 169:42]
  assign _T_429 = _T_123 & _T_428; // @[Parameters.scala 168:56]
  assign _T_431 = io_in_a_bits_size <= 4'h8; // @[Parameters.scala 90:42]
  assign _T_439 = _T_431 & _T_162; // @[Parameters.scala 168:56]
  assign _T_448 = _T_327 | _T_429; // @[Parameters.scala 170:30]
  assign _T_449 = _T_448 | _T_439; // @[Parameters.scala 170:30]
  assign _T_452 = _T_449 | reset; // @[Monitor.scala 81:14]
  assign _T_468 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 88:25]
  assign _T_542 = io_in_a_bits_mask & ~_T_100; // @[Monitor.scala 93:28]
  assign _T_543 = _T_542 == 8'h0; // @[Monitor.scala 93:37]
  assign _T_545 = _T_543 | reset; // @[Monitor.scala 93:14]
  assign _T_547 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 96:25]
  assign _T_549 = io_in_a_bits_size <= 4'h3; // @[Parameters.scala 90:42]
  assign _T_575 = _T_549 & _T_165; // @[Parameters.scala 168:56]
  assign _T_598 = _T_575 | reset; // @[Monitor.scala 97:14]
  assign _T_606 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 139:33]
  assign _T_608 = _T_606 | reset; // @[Monitor.scala 100:14]
  assign _T_614 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 104:25]
  assign _T_673 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 146:30]
  assign _T_675 = _T_673 | reset; // @[Monitor.scala 108:14]
  assign _T_681 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 112:25]
  assign _T_732 = _T_327 | reset; // @[Monitor.scala 113:14]
  assign _T_748 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 43:24]
  assign _T_750 = _T_748 | reset; // @[Monitor.scala 268:12]
  assign _T_762 = ~io_in_d_bits_source | io_in_d_bits_source; // @[Parameters.scala 280:46]
  assign _T_764 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 275:25]
  assign _T_766 = _T_762 | reset; // @[Monitor.scala 276:14]
  assign _T_768 = io_in_d_bits_size >= 4'h3; // @[Monitor.scala 277:27]
  assign _T_770 = _T_768 | reset; // @[Monitor.scala 277:14]
  assign _T_772 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 278:28]
  assign _T_774 = _T_772 | reset; // @[Monitor.scala 278:14]
  assign _T_778 = ~io_in_d_bits_corrupt | reset; // @[Monitor.scala 279:14]
  assign _T_782 = ~io_in_d_bits_denied | reset; // @[Monitor.scala 280:14]
  assign _T_784 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 283:25]
  assign _T_795 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 103:26]
  assign _T_797 = _T_795 | reset; // @[Monitor.scala 287:14]
  assign _T_799 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 288:28]
  assign _T_801 = _T_799 | reset; // @[Monitor.scala 288:14]
  assign _T_812 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 293:25]
  assign _T_832 = ~io_in_d_bits_denied | io_in_d_bits_corrupt; // @[Monitor.scala 299:30]
  assign _T_834 = _T_832 | reset; // @[Monitor.scala 299:14]
  assign _T_841 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 303:25]
  assign _T_858 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 311:25]
  assign _T_876 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 319:25]
  assign _T_893 = io_in_b_bits_opcode <= 3'h6; // @[Bundles.scala 41:24]
  assign _T_895 = _T_893 | reset; // @[Monitor.scala 122:12]
  assign _T_900 = {1'b0,$signed(io_in_b_bits_address)}; // @[Parameters.scala 121:49]
  assign _T_917 = io_in_b_bits_address ^ 32'h3000; // @[Parameters.scala 121:31]
  assign _T_918 = {1'b0,$signed(_T_917)}; // @[Parameters.scala 121:49]
  assign _T_920 = $signed(_T_918) & -33'sh1000; // @[Parameters.scala 121:52]
  assign _T_921 = $signed(_T_920) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_922 = io_in_b_bits_address ^ 32'hc000000; // @[Parameters.scala 121:31]
  assign _T_923 = {1'b0,$signed(_T_922)}; // @[Parameters.scala 121:49]
  assign _T_925 = $signed(_T_923) & -33'sh4000000; // @[Parameters.scala 121:52]
  assign _T_926 = $signed(_T_925) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_927 = io_in_b_bits_address ^ 32'h2000000; // @[Parameters.scala 121:31]
  assign _T_928 = {1'b0,$signed(_T_927)}; // @[Parameters.scala 121:49]
  assign _T_930 = $signed(_T_928) & -33'sh10000; // @[Parameters.scala 121:52]
  assign _T_931 = $signed(_T_930) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_935 = $signed(_T_900) & -33'sh1000; // @[Parameters.scala 121:52]
  assign _T_936 = $signed(_T_935) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_937 = io_in_b_bits_address ^ 32'h10000; // @[Parameters.scala 121:31]
  assign _T_938 = {1'b0,$signed(_T_937)}; // @[Parameters.scala 121:49]
  assign _T_940 = $signed(_T_938) & -33'sh10000; // @[Parameters.scala 121:52]
  assign _T_941 = $signed(_T_940) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_942 = io_in_b_bits_address ^ 32'h80000000; // @[Parameters.scala 121:31]
  assign _T_943 = {1'b0,$signed(_T_942)}; // @[Parameters.scala 121:49]
  assign _T_945 = $signed(_T_943) & -33'sh10000000; // @[Parameters.scala 121:52]
  assign _T_946 = $signed(_T_945) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_947 = io_in_b_bits_address ^ 32'h60000000; // @[Parameters.scala 121:31]
  assign _T_948 = {1'b0,$signed(_T_947)}; // @[Parameters.scala 121:49]
  assign _T_950 = $signed(_T_948) & -33'sh20000000; // @[Parameters.scala 121:52]
  assign _T_951 = $signed(_T_950) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_965 = _T_921 | _T_926; // @[Parameters.scala 155:64]
  assign _T_966 = _T_965 | _T_931; // @[Parameters.scala 155:64]
  assign _T_967 = _T_966 | _T_936; // @[Parameters.scala 155:64]
  assign _T_968 = _T_967 | _T_941; // @[Parameters.scala 155:64]
  assign _T_969 = _T_968 | _T_946; // @[Parameters.scala 155:64]
  assign _T_970 = _T_969 | _T_951; // @[Parameters.scala 155:64]
  assign _T_972 = 27'hfff << io_in_b_bits_size; // @[package.scala 185:77]
  assign _GEN_34 = {{20'd0}, ~_T_972[11:0]}; // @[Edges.scala 21:16]
  assign _T_975 = io_in_b_bits_address & _GEN_34; // @[Edges.scala 21:16]
  assign _T_976 = _T_975 == 32'h0; // @[Edges.scala 21:24]
  assign _T_979 = 4'h1 << io_in_b_bits_size[1:0]; // @[OneHot.scala 52:12]
  assign _T_981 = _T_979[2:0] | 3'h1; // @[Misc.scala 206:81]
  assign _T_982 = io_in_b_bits_size >= 4'h3; // @[Misc.scala 210:21]
  assign _T_987 = _T_981[2] & ~io_in_b_bits_address[2]; // @[Misc.scala 219:38]
  assign _T_988 = _T_982 | _T_987; // @[Misc.scala 219:29]
  assign _T_990 = _T_981[2] & io_in_b_bits_address[2]; // @[Misc.scala 219:38]
  assign _T_991 = _T_982 | _T_990; // @[Misc.scala 219:29]
  assign _T_995 = ~io_in_b_bits_address[2] & ~io_in_b_bits_address[1]; // @[Misc.scala 218:27]
  assign _T_996 = _T_981[1] & _T_995; // @[Misc.scala 219:38]
  assign _T_997 = _T_988 | _T_996; // @[Misc.scala 219:29]
  assign _T_998 = ~io_in_b_bits_address[2] & io_in_b_bits_address[1]; // @[Misc.scala 218:27]
  assign _T_999 = _T_981[1] & _T_998; // @[Misc.scala 219:38]
  assign _T_1000 = _T_988 | _T_999; // @[Misc.scala 219:29]
  assign _T_1001 = io_in_b_bits_address[2] & ~io_in_b_bits_address[1]; // @[Misc.scala 218:27]
  assign _T_1002 = _T_981[1] & _T_1001; // @[Misc.scala 219:38]
  assign _T_1003 = _T_991 | _T_1002; // @[Misc.scala 219:29]
  assign _T_1004 = io_in_b_bits_address[2] & io_in_b_bits_address[1]; // @[Misc.scala 218:27]
  assign _T_1005 = _T_981[1] & _T_1004; // @[Misc.scala 219:38]
  assign _T_1006 = _T_991 | _T_1005; // @[Misc.scala 219:29]
  assign _T_1010 = _T_995 & ~io_in_b_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_1011 = _T_981[0] & _T_1010; // @[Misc.scala 219:38]
  assign _T_1012 = _T_997 | _T_1011; // @[Misc.scala 219:29]
  assign _T_1013 = _T_995 & io_in_b_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_1014 = _T_981[0] & _T_1013; // @[Misc.scala 219:38]
  assign _T_1015 = _T_997 | _T_1014; // @[Misc.scala 219:29]
  assign _T_1016 = _T_998 & ~io_in_b_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_1017 = _T_981[0] & _T_1016; // @[Misc.scala 219:38]
  assign _T_1018 = _T_1000 | _T_1017; // @[Misc.scala 219:29]
  assign _T_1019 = _T_998 & io_in_b_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_1020 = _T_981[0] & _T_1019; // @[Misc.scala 219:38]
  assign _T_1021 = _T_1000 | _T_1020; // @[Misc.scala 219:29]
  assign _T_1022 = _T_1001 & ~io_in_b_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_1023 = _T_981[0] & _T_1022; // @[Misc.scala 219:38]
  assign _T_1024 = _T_1003 | _T_1023; // @[Misc.scala 219:29]
  assign _T_1025 = _T_1001 & io_in_b_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_1026 = _T_981[0] & _T_1025; // @[Misc.scala 219:38]
  assign _T_1027 = _T_1003 | _T_1026; // @[Misc.scala 219:29]
  assign _T_1028 = _T_1004 & ~io_in_b_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_1029 = _T_981[0] & _T_1028; // @[Misc.scala 219:38]
  assign _T_1030 = _T_1006 | _T_1029; // @[Misc.scala 219:29]
  assign _T_1031 = _T_1004 & io_in_b_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_1032 = _T_981[0] & _T_1031; // @[Misc.scala 219:38]
  assign _T_1033 = _T_1006 | _T_1032; // @[Misc.scala 219:29]
  assign _T_1040 = {_T_1033,_T_1030,_T_1027,_T_1024,_T_1021,_T_1018,_T_1015,_T_1012}; // @[Cat.scala 30:58]
  assign _T_1057 = io_in_b_bits_source == io_in_b_bits_source; // @[Monitor.scala 130:117]
  assign _T_1058 = io_in_b_bits_opcode == 3'h6; // @[Monitor.scala 132:25]
  assign _T_1069 = 4'h6 == io_in_b_bits_size; // @[Parameters.scala 89:48]
  assign _T_1071 = ~io_in_b_bits_source & _T_1069; // @[Mux.scala 19:72]
  assign _T_1077 = _T_1071 | reset; // @[Monitor.scala 133:14]
  assign _T_1080 = _T_970 | reset; // @[Monitor.scala 134:14]
  assign _T_1083 = _T_1057 | reset; // @[Monitor.scala 135:14]
  assign _T_1086 = _T_976 | reset; // @[Monitor.scala 136:14]
  assign _T_1088 = io_in_b_bits_param <= 2'h2; // @[Bundles.scala 103:26]
  assign _T_1090 = _T_1088 | reset; // @[Monitor.scala 137:14]
  assign _T_1092 = io_in_b_bits_mask == _T_1040; // @[Monitor.scala 138:27]
  assign _T_1094 = _T_1092 | reset; // @[Monitor.scala 138:14]
  assign _T_1098 = ~io_in_b_bits_corrupt | reset; // @[Monitor.scala 139:14]
  assign _T_1100 = io_in_b_bits_opcode == 3'h4; // @[Monitor.scala 142:25]
  assign _T_1113 = io_in_b_bits_param == 2'h0; // @[Monitor.scala 147:28]
  assign _T_1115 = _T_1113 | reset; // @[Monitor.scala 147:14]
  assign _T_1125 = io_in_b_bits_opcode == 3'h0; // @[Monitor.scala 152:25]
  assign _T_1146 = io_in_b_bits_opcode == 3'h1; // @[Monitor.scala 161:25]
  assign _T_1164 = io_in_b_bits_mask & ~_T_1040; // @[Monitor.scala 167:28]
  assign _T_1165 = _T_1164 == 8'h0; // @[Monitor.scala 167:37]
  assign _T_1167 = _T_1165 | reset; // @[Monitor.scala 167:14]
  assign _T_1169 = io_in_b_bits_opcode == 3'h2; // @[Monitor.scala 170:25]
  assign _T_1190 = io_in_b_bits_opcode == 3'h3; // @[Monitor.scala 179:25]
  assign _T_1211 = io_in_b_bits_opcode == 3'h5; // @[Monitor.scala 188:25]
  assign _T_1246 = ~io_in_c_bits_source | io_in_c_bits_source; // @[Parameters.scala 280:46]
  assign _T_1248 = 27'hfff << io_in_c_bits_size; // @[package.scala 185:77]
  assign _GEN_35 = {{20'd0}, ~_T_1248[11:0]}; // @[Edges.scala 21:16]
  assign _T_1251 = io_in_c_bits_address & _GEN_35; // @[Edges.scala 21:16]
  assign _T_1252 = _T_1251 == 32'h0; // @[Edges.scala 21:24]
  assign _T_1253 = io_in_c_bits_address ^ 32'h3000; // @[Parameters.scala 121:31]
  assign _T_1254 = {1'b0,$signed(_T_1253)}; // @[Parameters.scala 121:49]
  assign _T_1256 = $signed(_T_1254) & -33'sh1000; // @[Parameters.scala 121:52]
  assign _T_1257 = $signed(_T_1256) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_1258 = io_in_c_bits_address ^ 32'hc000000; // @[Parameters.scala 121:31]
  assign _T_1259 = {1'b0,$signed(_T_1258)}; // @[Parameters.scala 121:49]
  assign _T_1261 = $signed(_T_1259) & -33'sh4000000; // @[Parameters.scala 121:52]
  assign _T_1262 = $signed(_T_1261) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_1263 = io_in_c_bits_address ^ 32'h2000000; // @[Parameters.scala 121:31]
  assign _T_1264 = {1'b0,$signed(_T_1263)}; // @[Parameters.scala 121:49]
  assign _T_1266 = $signed(_T_1264) & -33'sh10000; // @[Parameters.scala 121:52]
  assign _T_1267 = $signed(_T_1266) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_1269 = {1'b0,$signed(io_in_c_bits_address)}; // @[Parameters.scala 121:49]
  assign _T_1271 = $signed(_T_1269) & -33'sh1000; // @[Parameters.scala 121:52]
  assign _T_1272 = $signed(_T_1271) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_1273 = io_in_c_bits_address ^ 32'h10000; // @[Parameters.scala 121:31]
  assign _T_1274 = {1'b0,$signed(_T_1273)}; // @[Parameters.scala 121:49]
  assign _T_1276 = $signed(_T_1274) & -33'sh10000; // @[Parameters.scala 121:52]
  assign _T_1277 = $signed(_T_1276) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_1278 = io_in_c_bits_address ^ 32'h80000000; // @[Parameters.scala 121:31]
  assign _T_1279 = {1'b0,$signed(_T_1278)}; // @[Parameters.scala 121:49]
  assign _T_1281 = $signed(_T_1279) & -33'sh10000000; // @[Parameters.scala 121:52]
  assign _T_1282 = $signed(_T_1281) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_1283 = io_in_c_bits_address ^ 32'h60000000; // @[Parameters.scala 121:31]
  assign _T_1284 = {1'b0,$signed(_T_1283)}; // @[Parameters.scala 121:49]
  assign _T_1286 = $signed(_T_1284) & -33'sh20000000; // @[Parameters.scala 121:52]
  assign _T_1287 = $signed(_T_1286) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_1301 = _T_1257 | _T_1262; // @[Parameters.scala 155:64]
  assign _T_1302 = _T_1301 | _T_1267; // @[Parameters.scala 155:64]
  assign _T_1303 = _T_1302 | _T_1272; // @[Parameters.scala 155:64]
  assign _T_1304 = _T_1303 | _T_1277; // @[Parameters.scala 155:64]
  assign _T_1305 = _T_1304 | _T_1282; // @[Parameters.scala 155:64]
  assign _T_1306 = _T_1305 | _T_1287; // @[Parameters.scala 155:64]
  assign _T_1327 = io_in_c_bits_opcode == 3'h4; // @[Monitor.scala 207:25]
  assign _T_1329 = _T_1306 | reset; // @[Monitor.scala 208:14]
  assign _T_1332 = _T_1246 | reset; // @[Monitor.scala 209:14]
  assign _T_1334 = io_in_c_bits_size >= 4'h3; // @[Monitor.scala 210:27]
  assign _T_1336 = _T_1334 | reset; // @[Monitor.scala 210:14]
  assign _T_1339 = _T_1252 | reset; // @[Monitor.scala 211:14]
  assign _T_1341 = io_in_c_bits_param <= 3'h5; // @[Bundles.scala 121:29]
  assign _T_1343 = _T_1341 | reset; // @[Monitor.scala 212:14]
  assign _T_1349 = io_in_c_bits_opcode == 3'h5; // @[Monitor.scala 216:25]
  assign _T_1367 = io_in_c_bits_opcode == 3'h6; // @[Monitor.scala 224:25]
  assign _T_1369 = io_in_c_bits_size <= 4'h6; // @[Parameters.scala 90:42]
  assign _T_1377 = _T_1369 & _T_1282; // @[Parameters.scala 168:56]
  assign _T_1418 = _T_1377 | reset; // @[Monitor.scala 225:14]
  assign _T_1430 = 4'h6 == io_in_c_bits_size; // @[Parameters.scala 89:48]
  assign _T_1432 = ~io_in_c_bits_source & _T_1430; // @[Mux.scala 19:72]
  assign _T_1438 = _T_1432 | reset; // @[Monitor.scala 226:14]
  assign _T_1450 = io_in_c_bits_param <= 3'h2; // @[Bundles.scala 115:29]
  assign _T_1452 = _T_1450 | reset; // @[Monitor.scala 230:14]
  assign _T_1458 = io_in_c_bits_opcode == 3'h7; // @[Monitor.scala 234:25]
  assign _T_1545 = io_in_c_bits_opcode == 3'h0; // @[Monitor.scala 243:25]
  assign _T_1555 = io_in_c_bits_param == 3'h0; // @[Monitor.scala 247:28]
  assign _T_1557 = _T_1555 | reset; // @[Monitor.scala 247:14]
  assign _T_1563 = io_in_c_bits_opcode == 3'h1; // @[Monitor.scala 251:25]
  assign _T_1577 = io_in_c_bits_opcode == 3'h2; // @[Monitor.scala 258:25]
  assign _T_1599 = io_in_a_ready & io_in_a_valid; // @[Bundles.scala 277:22]
  assign _T_1604 = ~_T_32[11:3]; // @[Edges.scala 220:59]
  assign _T_1612 = _T_1609 - 9'h1; // @[Edges.scala 230:28]
  assign _T_1613 = _T_1609 == 9'h0; // @[Edges.scala 231:25]
  assign _T_1632 = io_in_a_valid & ~_T_1613; // @[Monitor.scala 354:19]
  assign _T_1633 = io_in_a_bits_opcode == _T_1622; // @[Monitor.scala 355:29]
  assign _T_1635 = _T_1633 | reset; // @[Monitor.scala 355:14]
  assign _T_1637 = io_in_a_bits_param == _T_1624; // @[Monitor.scala 356:29]
  assign _T_1639 = _T_1637 | reset; // @[Monitor.scala 356:14]
  assign _T_1641 = io_in_a_bits_size == _T_1626; // @[Monitor.scala 357:29]
  assign _T_1643 = _T_1641 | reset; // @[Monitor.scala 357:14]
  assign _T_1645 = io_in_a_bits_source == _T_1628; // @[Monitor.scala 358:29]
  assign _T_1647 = _T_1645 | reset; // @[Monitor.scala 358:14]
  assign _T_1649 = io_in_a_bits_address == _T_1630; // @[Monitor.scala 359:29]
  assign _T_1651 = _T_1649 | reset; // @[Monitor.scala 359:14]
  assign _T_1654 = _T_1599 & _T_1613; // @[Monitor.scala 361:20]
  assign _T_1655 = io_in_d_ready & io_in_d_valid; // @[Bundles.scala 277:22]
  assign _T_1657 = 27'hfff << io_in_d_bits_size; // @[package.scala 185:77]
  assign _T_1660 = ~_T_1657[11:3]; // @[Edges.scala 220:59]
  assign _T_1667 = _T_1664 - 9'h1; // @[Edges.scala 230:28]
  assign _T_1668 = _T_1664 == 9'h0; // @[Edges.scala 231:25]
  assign _T_1689 = io_in_d_valid & ~_T_1668; // @[Monitor.scala 424:19]
  assign _T_1690 = io_in_d_bits_opcode == _T_1677; // @[Monitor.scala 425:29]
  assign _T_1692 = _T_1690 | reset; // @[Monitor.scala 425:14]
  assign _T_1694 = io_in_d_bits_param == _T_1679; // @[Monitor.scala 426:29]
  assign _T_1696 = _T_1694 | reset; // @[Monitor.scala 426:14]
  assign _T_1698 = io_in_d_bits_size == _T_1681; // @[Monitor.scala 427:29]
  assign _T_1700 = _T_1698 | reset; // @[Monitor.scala 427:14]
  assign _T_1702 = io_in_d_bits_source == _T_1683; // @[Monitor.scala 428:29]
  assign _T_1704 = _T_1702 | reset; // @[Monitor.scala 428:14]
  assign _T_1706 = io_in_d_bits_sink == _T_1685; // @[Monitor.scala 429:29]
  assign _T_1708 = _T_1706 | reset; // @[Monitor.scala 429:14]
  assign _T_1710 = io_in_d_bits_denied == _T_1687; // @[Monitor.scala 430:29]
  assign _T_1712 = _T_1710 | reset; // @[Monitor.scala 430:14]
  assign _T_1715 = _T_1655 & _T_1668; // @[Monitor.scala 432:20]
  assign _T_1716 = io_in_b_ready & io_in_b_valid; // @[Bundles.scala 277:22]
  assign _T_1729 = _T_1726 - 9'h1; // @[Edges.scala 230:28]
  assign _T_1730 = _T_1726 == 9'h0; // @[Edges.scala 231:25]
  assign _T_1749 = io_in_b_valid & ~_T_1730; // @[Monitor.scala 377:19]
  assign _T_1750 = io_in_b_bits_opcode == _T_1739; // @[Monitor.scala 378:29]
  assign _T_1752 = _T_1750 | reset; // @[Monitor.scala 378:14]
  assign _T_1754 = io_in_b_bits_param == _T_1741; // @[Monitor.scala 379:29]
  assign _T_1756 = _T_1754 | reset; // @[Monitor.scala 379:14]
  assign _T_1758 = io_in_b_bits_size == _T_1743; // @[Monitor.scala 380:29]
  assign _T_1760 = _T_1758 | reset; // @[Monitor.scala 380:14]
  assign _T_1762 = io_in_b_bits_source == _T_1745; // @[Monitor.scala 381:29]
  assign _T_1764 = _T_1762 | reset; // @[Monitor.scala 381:14]
  assign _T_1766 = io_in_b_bits_address == _T_1747; // @[Monitor.scala 382:29]
  assign _T_1768 = _T_1766 | reset; // @[Monitor.scala 382:14]
  assign _T_1771 = _T_1716 & _T_1730; // @[Monitor.scala 384:20]
  assign _T_1772 = io_in_c_ready & io_in_c_valid; // @[Bundles.scala 277:22]
  assign _T_1777 = ~_T_1248[11:3]; // @[Edges.scala 220:59]
  assign _T_1784 = _T_1781 - 9'h1; // @[Edges.scala 230:28]
  assign _T_1785 = _T_1781 == 9'h0; // @[Edges.scala 231:25]
  assign _T_1804 = io_in_c_valid & ~_T_1785; // @[Monitor.scala 400:19]
  assign _T_1805 = io_in_c_bits_opcode == _T_1794; // @[Monitor.scala 401:29]
  assign _T_1807 = _T_1805 | reset; // @[Monitor.scala 401:14]
  assign _T_1809 = io_in_c_bits_param == _T_1796; // @[Monitor.scala 402:29]
  assign _T_1811 = _T_1809 | reset; // @[Monitor.scala 402:14]
  assign _T_1813 = io_in_c_bits_size == _T_1798; // @[Monitor.scala 403:29]
  assign _T_1815 = _T_1813 | reset; // @[Monitor.scala 403:14]
  assign _T_1817 = io_in_c_bits_source == _T_1800; // @[Monitor.scala 404:29]
  assign _T_1819 = _T_1817 | reset; // @[Monitor.scala 404:14]
  assign _T_1821 = io_in_c_bits_address == _T_1802; // @[Monitor.scala 405:29]
  assign _T_1823 = _T_1821 | reset; // @[Monitor.scala 405:14]
  assign _T_1826 = _T_1772 & _T_1785; // @[Monitor.scala 407:20]
  assign _T_1842 = _T_1839 - 9'h1; // @[Edges.scala 230:28]
  assign _T_1843 = _T_1839 == 9'h0; // @[Edges.scala 231:25]
  assign _T_1863 = _T_1860 - 9'h1; // @[Edges.scala 230:28]
  assign _T_1864 = _T_1860 == 9'h0; // @[Edges.scala 231:25]
  assign _T_1875 = _T_1599 & _T_1843; // @[Monitor.scala 458:27]
  assign _T_1877 = 2'h1 << io_in_a_bits_source; // @[OneHot.scala 45:35]
  assign _T_1878 = _T_1828 >> io_in_a_bits_source; // @[Monitor.scala 460:23]
  assign _T_1882 = ~_T_1878[0] | reset; // @[Monitor.scala 460:13]
  assign _GEN_27 = _T_1875 ? _T_1877 : 2'h0; // @[Monitor.scala 458:72]
  assign _T_1888 = _T_1655 & _T_1864; // @[Monitor.scala 465:27]
  assign _T_1891 = _T_1888 & ~_T_764; // @[Monitor.scala 465:72]
  assign _T_1892 = 2'h1 << io_in_d_bits_source; // @[OneHot.scala 45:35]
  assign _T_1893 = _GEN_27 | _T_1828; // @[Monitor.scala 467:21]
  assign _T_1894 = _T_1893 >> io_in_d_bits_source; // @[Monitor.scala 467:32]
  assign _T_1897 = _T_1894[0] | reset; // @[Monitor.scala 467:13]
  assign _GEN_28 = _T_1891 ? _T_1892 : 2'h0; // @[Monitor.scala 465:91]
  assign _T_1899 = _GEN_27 != _GEN_28; // @[Monitor.scala 471:20]
  assign _T_1900 = _GEN_27 != 2'h0; // @[Monitor.scala 471:40]
  assign _T_1902 = _T_1899 | ~_T_1900; // @[Monitor.scala 471:30]
  assign _T_1904 = _T_1902 | reset; // @[Monitor.scala 471:13]
  assign _T_1906 = _T_1828 | _GEN_27; // @[Monitor.scala 474:27]
  assign _T_1908 = _T_1906 & ~_GEN_28; // @[Monitor.scala 474:36]
  assign _T_1939 = _T_1936 - 9'h1; // @[Edges.scala 230:28]
  assign _T_1940 = _T_1936 == 9'h0; // @[Edges.scala 231:25]
  assign _T_1951 = _T_1655 & _T_1940; // @[Monitor.scala 492:27]
  assign _T_1955 = io_in_d_bits_opcode[2] & ~io_in_d_bits_opcode[1]; // @[Edges.scala 71:40]
  assign _T_1956 = _T_1951 & _T_1955; // @[Monitor.scala 492:38]
  assign _T_1957 = 4'h1 << io_in_d_bits_sink; // @[OneHot.scala 45:35]
  assign _T_1958 = _T_1926 >> io_in_d_bits_sink; // @[Monitor.scala 494:23]
  assign _T_1962 = ~_T_1958[0] | reset; // @[Monitor.scala 494:13]
  assign _GEN_31 = _T_1956 ? _T_1957 : 4'h0; // @[Monitor.scala 492:72]
  assign _T_1966 = io_in_e_ready & io_in_e_valid; // @[Bundles.scala 277:22]
  assign _T_1969 = 4'h1 << io_in_e_bits_sink; // @[OneHot.scala 45:35]
  assign _T_1970 = _GEN_31 | _T_1926; // @[Monitor.scala 500:21]
  assign _T_1971 = _T_1970 >> io_in_e_bits_sink; // @[Monitor.scala 500:32]
  assign _T_1974 = _T_1971[0] | reset; // @[Monitor.scala 500:13]
  assign _GEN_32 = _T_1966 ? _T_1969 : 4'h0; // @[Monitor.scala 498:73]
  assign _T_1976 = _T_1926 | _GEN_31; // @[Monitor.scala 505:27]
  assign _T_1978 = _T_1976 & ~_GEN_32; // @[Monitor.scala 505:36]
  assign _GEN_36 = io_in_a_valid & _T_121; // @[Monitor.scala 49:14]
  assign _GEN_50 = io_in_a_valid & _T_217; // @[Monitor.scala 60:14]
  assign _GEN_66 = io_in_a_valid & _T_317; // @[Monitor.scala 72:14]
  assign _GEN_76 = io_in_a_valid & _T_391; // @[Monitor.scala 81:14]
  assign _GEN_86 = io_in_a_valid & _T_468; // @[Monitor.scala 89:14]
  assign _GEN_96 = io_in_a_valid & _T_547; // @[Monitor.scala 97:14]
  assign _GEN_106 = io_in_a_valid & _T_614; // @[Monitor.scala 105:14]
  assign _GEN_116 = io_in_a_valid & _T_681; // @[Monitor.scala 113:14]
  assign _GEN_124 = io_in_d_valid & _T_764; // @[Monitor.scala 276:14]
  assign _GEN_134 = io_in_d_valid & _T_784; // @[Monitor.scala 284:14]
  assign _GEN_144 = io_in_d_valid & _T_812; // @[Monitor.scala 294:14]
  assign _GEN_154 = io_in_d_valid & _T_841; // @[Monitor.scala 304:14]
  assign _GEN_160 = io_in_d_valid & _T_858; // @[Monitor.scala 312:14]
  assign _GEN_166 = io_in_d_valid & _T_876; // @[Monitor.scala 320:14]
  assign _GEN_172 = io_in_b_valid & _T_1058; // @[Monitor.scala 133:14]
  assign _GEN_186 = io_in_b_valid & _T_1100; // @[Monitor.scala 143:14]
  assign _GEN_200 = io_in_b_valid & _T_1125; // @[Monitor.scala 153:14]
  assign _GEN_212 = io_in_b_valid & _T_1146; // @[Monitor.scala 162:14]
  assign _GEN_224 = io_in_b_valid & _T_1169; // @[Monitor.scala 171:14]
  assign _GEN_234 = io_in_b_valid & _T_1190; // @[Monitor.scala 180:14]
  assign _GEN_244 = io_in_b_valid & _T_1211; // @[Monitor.scala 189:14]
  assign _GEN_256 = io_in_c_valid & _T_1327; // @[Monitor.scala 208:14]
  assign _GEN_266 = io_in_c_valid & _T_1349; // @[Monitor.scala 217:14]
  assign _GEN_276 = io_in_c_valid & _T_1367; // @[Monitor.scala 225:14]
  assign _GEN_288 = io_in_c_valid & _T_1458; // @[Monitor.scala 235:14]
  assign _GEN_300 = io_in_c_valid & _T_1545; // @[Monitor.scala 244:14]
  assign _GEN_308 = io_in_c_valid & _T_1563; // @[Monitor.scala 252:14]
  assign _GEN_316 = io_in_c_valid & _T_1577; // @[Monitor.scala 259:14]
  assign TLMonitor_64_covSum = 30'h0;
  assign io_covSum = TLMonitor_64_covSum;
  assign stopEn0 = _GEN_36 & ~_T_172;
  assign stopEn1 = _GEN_36 & ~_T_192;
  assign stopEn2 = _GEN_36 & ~_T_195;
  assign stopEn3 = _GEN_36 & ~_T_199;
  assign stopEn4 = _GEN_36 & ~_T_202;
  assign stopEn5 = _GEN_36 & ~_T_206;
  assign stopEn6 = _GEN_36 & ~_T_211;
  assign stopEn7 = _GEN_50 & ~_T_172;
  assign stopEn8 = _GEN_50 & ~_T_192;
  assign stopEn9 = _GEN_50 & ~_T_195;
  assign stopEn10 = _GEN_50 & ~_T_199;
  assign stopEn11 = _GEN_50 & ~_T_202;
  assign stopEn12 = _GEN_50 & ~_T_206;
  assign stopEn13 = _GEN_50 & ~_T_306;
  assign stopEn14 = _GEN_50 & ~_T_211;
  assign stopEn15 = _GEN_66 & ~_T_371;
  assign stopEn16 = _GEN_66 & ~_T_195;
  assign stopEn17 = _GEN_66 & ~_T_202;
  assign stopEn18 = _GEN_66 & ~_T_381;
  assign stopEn19 = _GEN_66 & ~_T_385;
  assign stopEn20 = _GEN_76 & ~_T_452;
  assign stopEn21 = _GEN_76 & ~_T_195;
  assign stopEn22 = _GEN_76 & ~_T_202;
  assign stopEn23 = _GEN_76 & ~_T_381;
  assign stopEn24 = _GEN_76 & ~_T_385;
  assign stopEn25 = _GEN_86 & ~_T_452;
  assign stopEn26 = _GEN_86 & ~_T_195;
  assign stopEn27 = _GEN_86 & ~_T_202;
  assign stopEn28 = _GEN_86 & ~_T_381;
  assign stopEn29 = _GEN_86 & ~_T_545;
  assign stopEn30 = _GEN_96 & ~_T_598;
  assign stopEn31 = _GEN_96 & ~_T_195;
  assign stopEn32 = _GEN_96 & ~_T_202;
  assign stopEn33 = _GEN_96 & ~_T_608;
  assign stopEn34 = _GEN_96 & ~_T_385;
  assign stopEn35 = _GEN_106 & ~_T_598;
  assign stopEn36 = _GEN_106 & ~_T_195;
  assign stopEn37 = _GEN_106 & ~_T_202;
  assign stopEn38 = _GEN_106 & ~_T_675;
  assign stopEn39 = _GEN_106 & ~_T_385;
  assign stopEn40 = _GEN_116 & ~_T_732;
  assign stopEn41 = _GEN_116 & ~_T_195;
  assign stopEn42 = _GEN_116 & ~_T_202;
  assign stopEn43 = _GEN_116 & ~_T_385;
  assign stopEn44 = io_in_d_valid & ~_T_750;
  assign stopEn45 = _GEN_124 & ~_T_766;
  assign stopEn46 = _GEN_124 & ~_T_770;
  assign stopEn47 = _GEN_124 & ~_T_774;
  assign stopEn48 = _GEN_124 & ~_T_778;
  assign stopEn49 = _GEN_124 & ~_T_782;
  assign stopEn50 = _GEN_134 & ~_T_766;
  assign stopEn51 = _GEN_134 & ~_T_770;
  assign stopEn52 = _GEN_134 & ~_T_797;
  assign stopEn53 = _GEN_134 & ~_T_801;
  assign stopEn54 = _GEN_134 & ~_T_778;
  assign stopEn55 = _GEN_144 & ~_T_766;
  assign stopEn56 = _GEN_144 & ~_T_770;
  assign stopEn57 = _GEN_144 & ~_T_797;
  assign stopEn58 = _GEN_144 & ~_T_801;
  assign stopEn59 = _GEN_144 & ~_T_834;
  assign stopEn60 = _GEN_154 & ~_T_766;
  assign stopEn61 = _GEN_154 & ~_T_774;
  assign stopEn62 = _GEN_154 & ~_T_778;
  assign stopEn63 = _GEN_160 & ~_T_766;
  assign stopEn64 = _GEN_160 & ~_T_774;
  assign stopEn65 = _GEN_160 & ~_T_834;
  assign stopEn66 = _GEN_166 & ~_T_766;
  assign stopEn67 = _GEN_166 & ~_T_774;
  assign stopEn68 = _GEN_166 & ~_T_778;
  assign stopEn69 = io_in_b_valid & ~_T_895;
  assign stopEn70 = _GEN_172 & ~_T_1077;
  assign stopEn71 = _GEN_172 & ~_T_1080;
  assign stopEn72 = _GEN_172 & ~_T_1083;
  assign stopEn73 = _GEN_172 & ~_T_1086;
  assign stopEn74 = _GEN_172 & ~_T_1090;
  assign stopEn75 = _GEN_172 & ~_T_1094;
  assign stopEn76 = _GEN_172 & ~_T_1098;
  assign stopEn77 = _GEN_186 & ~reset;
  assign stopEn78 = _GEN_186 & ~_T_1080;
  assign stopEn79 = _GEN_186 & ~_T_1083;
  assign stopEn80 = _GEN_186 & ~_T_1086;
  assign stopEn81 = _GEN_186 & ~_T_1115;
  assign stopEn82 = _GEN_186 & ~_T_1094;
  assign stopEn83 = _GEN_186 & ~_T_1098;
  assign stopEn84 = _GEN_200 & ~reset;
  assign stopEn85 = _GEN_200 & ~_T_1080;
  assign stopEn86 = _GEN_200 & ~_T_1083;
  assign stopEn87 = _GEN_200 & ~_T_1086;
  assign stopEn88 = _GEN_200 & ~_T_1115;
  assign stopEn89 = _GEN_200 & ~_T_1094;
  assign stopEn90 = _GEN_212 & ~reset;
  assign stopEn91 = _GEN_212 & ~_T_1080;
  assign stopEn92 = _GEN_212 & ~_T_1083;
  assign stopEn93 = _GEN_212 & ~_T_1086;
  assign stopEn94 = _GEN_212 & ~_T_1115;
  assign stopEn95 = _GEN_212 & ~_T_1167;
  assign stopEn96 = _GEN_224 & ~reset;
  assign stopEn97 = _GEN_224 & ~_T_1080;
  assign stopEn98 = _GEN_224 & ~_T_1083;
  assign stopEn99 = _GEN_224 & ~_T_1086;
  assign stopEn100 = _GEN_224 & ~_T_1094;
  assign stopEn101 = _GEN_234 & ~reset;
  assign stopEn102 = _GEN_234 & ~_T_1080;
  assign stopEn103 = _GEN_234 & ~_T_1083;
  assign stopEn104 = _GEN_234 & ~_T_1086;
  assign stopEn105 = _GEN_234 & ~_T_1094;
  assign stopEn106 = _GEN_244 & ~reset;
  assign stopEn107 = _GEN_244 & ~_T_1080;
  assign stopEn108 = _GEN_244 & ~_T_1083;
  assign stopEn109 = _GEN_244 & ~_T_1086;
  assign stopEn110 = _GEN_244 & ~_T_1094;
  assign stopEn111 = _GEN_244 & ~_T_1098;
  assign stopEn112 = _GEN_256 & ~_T_1329;
  assign stopEn113 = _GEN_256 & ~_T_1332;
  assign stopEn114 = _GEN_256 & ~_T_1336;
  assign stopEn115 = _GEN_256 & ~_T_1339;
  assign stopEn116 = _GEN_256 & ~_T_1343;
  assign stopEn117 = _GEN_266 & ~_T_1329;
  assign stopEn118 = _GEN_266 & ~_T_1332;
  assign stopEn119 = _GEN_266 & ~_T_1336;
  assign stopEn120 = _GEN_266 & ~_T_1339;
  assign stopEn121 = _GEN_266 & ~_T_1343;
  assign stopEn122 = _GEN_276 & ~_T_1418;
  assign stopEn123 = _GEN_276 & ~_T_1438;
  assign stopEn124 = _GEN_276 & ~_T_1332;
  assign stopEn125 = _GEN_276 & ~_T_1336;
  assign stopEn126 = _GEN_276 & ~_T_1339;
  assign stopEn127 = _GEN_276 & ~_T_1452;
  assign stopEn128 = _GEN_288 & ~_T_1418;
  assign stopEn129 = _GEN_288 & ~_T_1438;
  assign stopEn130 = _GEN_288 & ~_T_1332;
  assign stopEn131 = _GEN_288 & ~_T_1336;
  assign stopEn132 = _GEN_288 & ~_T_1339;
  assign stopEn133 = _GEN_288 & ~_T_1452;
  assign stopEn134 = _GEN_300 & ~_T_1329;
  assign stopEn135 = _GEN_300 & ~_T_1332;
  assign stopEn136 = _GEN_300 & ~_T_1339;
  assign stopEn137 = _GEN_300 & ~_T_1557;
  assign stopEn138 = _GEN_308 & ~_T_1329;
  assign stopEn139 = _GEN_308 & ~_T_1332;
  assign stopEn140 = _GEN_308 & ~_T_1339;
  assign stopEn141 = _GEN_308 & ~_T_1557;
  assign stopEn142 = _GEN_316 & ~_T_1329;
  assign stopEn143 = _GEN_316 & ~_T_1332;
  assign stopEn144 = _GEN_316 & ~_T_1339;
  assign stopEn145 = _GEN_316 & ~_T_1557;
  assign stopEn146 = _T_1632 & ~_T_1635;
  assign stopEn147 = _T_1632 & ~_T_1639;
  assign stopEn148 = _T_1632 & ~_T_1643;
  assign stopEn149 = _T_1632 & ~_T_1647;
  assign stopEn150 = _T_1632 & ~_T_1651;
  assign stopEn151 = _T_1689 & ~_T_1692;
  assign stopEn152 = _T_1689 & ~_T_1696;
  assign stopEn153 = _T_1689 & ~_T_1700;
  assign stopEn154 = _T_1689 & ~_T_1704;
  assign stopEn155 = _T_1689 & ~_T_1708;
  assign stopEn156 = _T_1689 & ~_T_1712;
  assign stopEn157 = _T_1749 & ~_T_1752;
  assign stopEn158 = _T_1749 & ~_T_1756;
  assign stopEn159 = _T_1749 & ~_T_1760;
  assign stopEn160 = _T_1749 & ~_T_1764;
  assign stopEn161 = _T_1749 & ~_T_1768;
  assign stopEn162 = _T_1804 & ~_T_1807;
  assign stopEn163 = _T_1804 & ~_T_1811;
  assign stopEn164 = _T_1804 & ~_T_1815;
  assign stopEn165 = _T_1804 & ~_T_1819;
  assign stopEn166 = _T_1804 & ~_T_1823;
  assign stopEn167 = _T_1875 & ~_T_1882;
  assign stopEn168 = _T_1891 & ~_T_1897;
  assign stopEn169 = ~_T_1904;
  assign stopEn170 = _T_1956 & ~_T_1962;
  assign stopEn171 = _T_1966 & ~_T_1974;
  assign TLMonitor_64_or63 = stopEn0 | stopEn1;
  assign TLMonitor_64_or130 = stopEn3 | stopEn4;
  assign TLMonitor_64_or64 = stopEn2 | TLMonitor_64_or130;
  assign TLMonitor_64_or31 = TLMonitor_64_or63 | TLMonitor_64_or64;
  assign TLMonitor_64_or65 = stopEn5 | stopEn6;
  assign TLMonitor_64_or134 = stopEn8 | stopEn9;
  assign TLMonitor_64_or66 = stopEn7 | TLMonitor_64_or134;
  assign TLMonitor_64_or32 = TLMonitor_64_or65 | TLMonitor_64_or66;
  assign TLMonitor_64_or15 = TLMonitor_64_or31 | TLMonitor_64_or32;
  assign TLMonitor_64_or67 = stopEn10 | stopEn11;
  assign TLMonitor_64_or138 = stopEn13 | stopEn14;
  assign TLMonitor_64_or68 = stopEn12 | TLMonitor_64_or138;
  assign TLMonitor_64_or33 = TLMonitor_64_or67 | TLMonitor_64_or68;
  assign TLMonitor_64_or140 = stopEn16 | stopEn17;
  assign TLMonitor_64_or69 = stopEn15 | TLMonitor_64_or140;
  assign TLMonitor_64_or142 = stopEn19 | stopEn20;
  assign TLMonitor_64_or70 = stopEn18 | TLMonitor_64_or142;
  assign TLMonitor_64_or34 = TLMonitor_64_or69 | TLMonitor_64_or70;
  assign TLMonitor_64_or16 = TLMonitor_64_or33 | TLMonitor_64_or34;
  assign TLMonitor_64_or7 = TLMonitor_64_or15 | TLMonitor_64_or16;
  assign TLMonitor_64_or71 = stopEn21 | stopEn22;
  assign TLMonitor_64_or146 = stopEn24 | stopEn25;
  assign TLMonitor_64_or72 = stopEn23 | TLMonitor_64_or146;
  assign TLMonitor_64_or35 = TLMonitor_64_or71 | TLMonitor_64_or72;
  assign TLMonitor_64_or148 = stopEn27 | stopEn28;
  assign TLMonitor_64_or73 = stopEn26 | TLMonitor_64_or148;
  assign TLMonitor_64_or150 = stopEn30 | stopEn31;
  assign TLMonitor_64_or74 = stopEn29 | TLMonitor_64_or150;
  assign TLMonitor_64_or36 = TLMonitor_64_or73 | TLMonitor_64_or74;
  assign TLMonitor_64_or17 = TLMonitor_64_or35 | TLMonitor_64_or36;
  assign TLMonitor_64_or75 = stopEn32 | stopEn33;
  assign TLMonitor_64_or154 = stopEn35 | stopEn36;
  assign TLMonitor_64_or76 = stopEn34 | TLMonitor_64_or154;
  assign TLMonitor_64_or37 = TLMonitor_64_or75 | TLMonitor_64_or76;
  assign TLMonitor_64_or156 = stopEn38 | stopEn39;
  assign TLMonitor_64_or77 = stopEn37 | TLMonitor_64_or156;
  assign TLMonitor_64_or158 = stopEn41 | stopEn42;
  assign TLMonitor_64_or78 = stopEn40 | TLMonitor_64_or158;
  assign TLMonitor_64_or38 = TLMonitor_64_or77 | TLMonitor_64_or78;
  assign TLMonitor_64_or18 = TLMonitor_64_or37 | TLMonitor_64_or38;
  assign TLMonitor_64_or8 = TLMonitor_64_or17 | TLMonitor_64_or18;
  assign TLMonitor_64_or3 = TLMonitor_64_or7 | TLMonitor_64_or8;
  assign TLMonitor_64_or79 = stopEn43 | stopEn44;
  assign TLMonitor_64_or162 = stopEn46 | stopEn47;
  assign TLMonitor_64_or80 = stopEn45 | TLMonitor_64_or162;
  assign TLMonitor_64_or39 = TLMonitor_64_or79 | TLMonitor_64_or80;
  assign TLMonitor_64_or81 = stopEn48 | stopEn49;
  assign TLMonitor_64_or166 = stopEn51 | stopEn52;
  assign TLMonitor_64_or82 = stopEn50 | TLMonitor_64_or166;
  assign TLMonitor_64_or40 = TLMonitor_64_or81 | TLMonitor_64_or82;
  assign TLMonitor_64_or19 = TLMonitor_64_or39 | TLMonitor_64_or40;
  assign TLMonitor_64_or83 = stopEn53 | stopEn54;
  assign TLMonitor_64_or170 = stopEn56 | stopEn57;
  assign TLMonitor_64_or84 = stopEn55 | TLMonitor_64_or170;
  assign TLMonitor_64_or41 = TLMonitor_64_or83 | TLMonitor_64_or84;
  assign TLMonitor_64_or172 = stopEn59 | stopEn60;
  assign TLMonitor_64_or85 = stopEn58 | TLMonitor_64_or172;
  assign TLMonitor_64_or174 = stopEn62 | stopEn63;
  assign TLMonitor_64_or86 = stopEn61 | TLMonitor_64_or174;
  assign TLMonitor_64_or42 = TLMonitor_64_or85 | TLMonitor_64_or86;
  assign TLMonitor_64_or20 = TLMonitor_64_or41 | TLMonitor_64_or42;
  assign TLMonitor_64_or9 = TLMonitor_64_or19 | TLMonitor_64_or20;
  assign TLMonitor_64_or87 = stopEn64 | stopEn65;
  assign TLMonitor_64_or178 = stopEn67 | stopEn68;
  assign TLMonitor_64_or88 = stopEn66 | TLMonitor_64_or178;
  assign TLMonitor_64_or43 = TLMonitor_64_or87 | TLMonitor_64_or88;
  assign TLMonitor_64_or180 = stopEn70 | stopEn71;
  assign TLMonitor_64_or89 = stopEn69 | TLMonitor_64_or180;
  assign TLMonitor_64_or182 = stopEn73 | stopEn74;
  assign TLMonitor_64_or90 = stopEn72 | TLMonitor_64_or182;
  assign TLMonitor_64_or44 = TLMonitor_64_or89 | TLMonitor_64_or90;
  assign TLMonitor_64_or21 = TLMonitor_64_or43 | TLMonitor_64_or44;
  assign TLMonitor_64_or91 = stopEn75 | stopEn76;
  assign TLMonitor_64_or186 = stopEn78 | stopEn79;
  assign TLMonitor_64_or92 = stopEn77 | TLMonitor_64_or186;
  assign TLMonitor_64_or45 = TLMonitor_64_or91 | TLMonitor_64_or92;
  assign TLMonitor_64_or188 = stopEn81 | stopEn82;
  assign TLMonitor_64_or93 = stopEn80 | TLMonitor_64_or188;
  assign TLMonitor_64_or190 = stopEn84 | stopEn85;
  assign TLMonitor_64_or94 = stopEn83 | TLMonitor_64_or190;
  assign TLMonitor_64_or46 = TLMonitor_64_or93 | TLMonitor_64_or94;
  assign TLMonitor_64_or22 = TLMonitor_64_or45 | TLMonitor_64_or46;
  assign TLMonitor_64_or10 = TLMonitor_64_or21 | TLMonitor_64_or22;
  assign TLMonitor_64_or4 = TLMonitor_64_or9 | TLMonitor_64_or10;
  assign TLMonitor_64_or1 = TLMonitor_64_or3 | TLMonitor_64_or4;
  assign TLMonitor_64_or95 = stopEn86 | stopEn87;
  assign TLMonitor_64_or194 = stopEn89 | stopEn90;
  assign TLMonitor_64_or96 = stopEn88 | TLMonitor_64_or194;
  assign TLMonitor_64_or47 = TLMonitor_64_or95 | TLMonitor_64_or96;
  assign TLMonitor_64_or97 = stopEn91 | stopEn92;
  assign TLMonitor_64_or198 = stopEn94 | stopEn95;
  assign TLMonitor_64_or98 = stopEn93 | TLMonitor_64_or198;
  assign TLMonitor_64_or48 = TLMonitor_64_or97 | TLMonitor_64_or98;
  assign TLMonitor_64_or23 = TLMonitor_64_or47 | TLMonitor_64_or48;
  assign TLMonitor_64_or99 = stopEn96 | stopEn97;
  assign TLMonitor_64_or202 = stopEn99 | stopEn100;
  assign TLMonitor_64_or100 = stopEn98 | TLMonitor_64_or202;
  assign TLMonitor_64_or49 = TLMonitor_64_or99 | TLMonitor_64_or100;
  assign TLMonitor_64_or204 = stopEn102 | stopEn103;
  assign TLMonitor_64_or101 = stopEn101 | TLMonitor_64_or204;
  assign TLMonitor_64_or206 = stopEn105 | stopEn106;
  assign TLMonitor_64_or102 = stopEn104 | TLMonitor_64_or206;
  assign TLMonitor_64_or50 = TLMonitor_64_or101 | TLMonitor_64_or102;
  assign TLMonitor_64_or24 = TLMonitor_64_or49 | TLMonitor_64_or50;
  assign TLMonitor_64_or11 = TLMonitor_64_or23 | TLMonitor_64_or24;
  assign TLMonitor_64_or103 = stopEn107 | stopEn108;
  assign TLMonitor_64_or210 = stopEn110 | stopEn111;
  assign TLMonitor_64_or104 = stopEn109 | TLMonitor_64_or210;
  assign TLMonitor_64_or51 = TLMonitor_64_or103 | TLMonitor_64_or104;
  assign TLMonitor_64_or212 = stopEn113 | stopEn114;
  assign TLMonitor_64_or105 = stopEn112 | TLMonitor_64_or212;
  assign TLMonitor_64_or214 = stopEn116 | stopEn117;
  assign TLMonitor_64_or106 = stopEn115 | TLMonitor_64_or214;
  assign TLMonitor_64_or52 = TLMonitor_64_or105 | TLMonitor_64_or106;
  assign TLMonitor_64_or25 = TLMonitor_64_or51 | TLMonitor_64_or52;
  assign TLMonitor_64_or107 = stopEn118 | stopEn119;
  assign TLMonitor_64_or218 = stopEn121 | stopEn122;
  assign TLMonitor_64_or108 = stopEn120 | TLMonitor_64_or218;
  assign TLMonitor_64_or53 = TLMonitor_64_or107 | TLMonitor_64_or108;
  assign TLMonitor_64_or220 = stopEn124 | stopEn125;
  assign TLMonitor_64_or109 = stopEn123 | TLMonitor_64_or220;
  assign TLMonitor_64_or222 = stopEn127 | stopEn128;
  assign TLMonitor_64_or110 = stopEn126 | TLMonitor_64_or222;
  assign TLMonitor_64_or54 = TLMonitor_64_or109 | TLMonitor_64_or110;
  assign TLMonitor_64_or26 = TLMonitor_64_or53 | TLMonitor_64_or54;
  assign TLMonitor_64_or12 = TLMonitor_64_or25 | TLMonitor_64_or26;
  assign TLMonitor_64_or5 = TLMonitor_64_or11 | TLMonitor_64_or12;
  assign TLMonitor_64_or111 = stopEn129 | stopEn130;
  assign TLMonitor_64_or226 = stopEn132 | stopEn133;
  assign TLMonitor_64_or112 = stopEn131 | TLMonitor_64_or226;
  assign TLMonitor_64_or55 = TLMonitor_64_or111 | TLMonitor_64_or112;
  assign TLMonitor_64_or113 = stopEn134 | stopEn135;
  assign TLMonitor_64_or230 = stopEn137 | stopEn138;
  assign TLMonitor_64_or114 = stopEn136 | TLMonitor_64_or230;
  assign TLMonitor_64_or56 = TLMonitor_64_or113 | TLMonitor_64_or114;
  assign TLMonitor_64_or27 = TLMonitor_64_or55 | TLMonitor_64_or56;
  assign TLMonitor_64_or115 = stopEn139 | stopEn140;
  assign TLMonitor_64_or234 = stopEn142 | stopEn143;
  assign TLMonitor_64_or116 = stopEn141 | TLMonitor_64_or234;
  assign TLMonitor_64_or57 = TLMonitor_64_or115 | TLMonitor_64_or116;
  assign TLMonitor_64_or236 = stopEn145 | stopEn146;
  assign TLMonitor_64_or117 = stopEn144 | TLMonitor_64_or236;
  assign TLMonitor_64_or238 = stopEn148 | stopEn149;
  assign TLMonitor_64_or118 = stopEn147 | TLMonitor_64_or238;
  assign TLMonitor_64_or58 = TLMonitor_64_or117 | TLMonitor_64_or118;
  assign TLMonitor_64_or28 = TLMonitor_64_or57 | TLMonitor_64_or58;
  assign TLMonitor_64_or13 = TLMonitor_64_or27 | TLMonitor_64_or28;
  assign TLMonitor_64_or119 = stopEn150 | stopEn151;
  assign TLMonitor_64_or242 = stopEn153 | stopEn154;
  assign TLMonitor_64_or120 = stopEn152 | TLMonitor_64_or242;
  assign TLMonitor_64_or59 = TLMonitor_64_or119 | TLMonitor_64_or120;
  assign TLMonitor_64_or244 = stopEn156 | stopEn157;
  assign TLMonitor_64_or121 = stopEn155 | TLMonitor_64_or244;
  assign TLMonitor_64_or246 = stopEn159 | stopEn160;
  assign TLMonitor_64_or122 = stopEn158 | TLMonitor_64_or246;
  assign TLMonitor_64_or60 = TLMonitor_64_or121 | TLMonitor_64_or122;
  assign TLMonitor_64_or29 = TLMonitor_64_or59 | TLMonitor_64_or60;
  assign TLMonitor_64_or123 = stopEn161 | stopEn162;
  assign TLMonitor_64_or250 = stopEn164 | stopEn165;
  assign TLMonitor_64_or124 = stopEn163 | TLMonitor_64_or250;
  assign TLMonitor_64_or61 = TLMonitor_64_or123 | TLMonitor_64_or124;
  assign TLMonitor_64_or252 = stopEn167 | stopEn168;
  assign TLMonitor_64_or125 = stopEn166 | TLMonitor_64_or252;
  assign TLMonitor_64_or254 = stopEn170 | stopEn171;
  assign TLMonitor_64_or126 = stopEn169 | TLMonitor_64_or254;
  assign TLMonitor_64_or62 = TLMonitor_64_or125 | TLMonitor_64_or126;
  assign TLMonitor_64_or30 = TLMonitor_64_or61 | TLMonitor_64_or62;
  assign TLMonitor_64_or14 = TLMonitor_64_or29 | TLMonitor_64_or30;
  assign TLMonitor_64_or6 = TLMonitor_64_or13 | TLMonitor_64_or14;
  assign TLMonitor_64_or2 = TLMonitor_64_or5 | TLMonitor_64_or6;
  assign TLMonitor_64_or0 = TLMonitor_64_or1 | TLMonitor_64_or2;
  assign metaAssert = TLMonitor_64_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1609 = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1622 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1624 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1626 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1628 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1630 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_1664 = _RAND_6[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_1677 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_1679 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_1681 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_1683 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_1685 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_1687 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_1726 = _RAND_13[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_1739 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_1741 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_1743 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_1745 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_1747 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_1781 = _RAND_19[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_1794 = _RAND_20[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_1796 = _RAND_21[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_1798 = _RAND_22[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_1800 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_1802 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_1828 = _RAND_25[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_1839 = _RAND_26[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_1860 = _RAND_27[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_1926 = _RAND_28[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_1936 = _RAND_29[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  TLMonitor_64_metaAssert = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      _T_1609 <= 9'h0;
    end else if (reset) begin
      _T_1609 <= 9'h0;
    end else if (_T_1599) begin
      if (_T_1613) begin
        if (~io_in_a_bits_opcode[2]) begin
          _T_1609 <= _T_1604;
        end else begin
          _T_1609 <= 9'h0;
        end
      end else begin
        _T_1609 <= _T_1612;
      end
    end
    if (metaReset) begin
      _T_1622 <= 3'h0;
    end else if (_T_1654) begin
      _T_1622 <= io_in_a_bits_opcode;
    end
    if (metaReset) begin
      _T_1624 <= 3'h0;
    end else if (_T_1654) begin
      _T_1624 <= io_in_a_bits_param;
    end
    if (metaReset) begin
      _T_1626 <= 4'h0;
    end else if (_T_1654) begin
      _T_1626 <= io_in_a_bits_size;
    end
    if (metaReset) begin
      _T_1628 <= 1'h0;
    end else if (_T_1654) begin
      _T_1628 <= io_in_a_bits_source;
    end
    if (metaReset) begin
      _T_1630 <= 32'h0;
    end else if (_T_1654) begin
      _T_1630 <= io_in_a_bits_address;
    end
    if (metaReset) begin
      _T_1664 <= 9'h0;
    end else if (reset) begin
      _T_1664 <= 9'h0;
    end else if (_T_1655) begin
      if (_T_1668) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1664 <= _T_1660;
        end else begin
          _T_1664 <= 9'h0;
        end
      end else begin
        _T_1664 <= _T_1667;
      end
    end
    if (metaReset) begin
      _T_1677 <= 3'h0;
    end else if (_T_1715) begin
      _T_1677 <= io_in_d_bits_opcode;
    end
    if (metaReset) begin
      _T_1679 <= 2'h0;
    end else if (_T_1715) begin
      _T_1679 <= io_in_d_bits_param;
    end
    if (metaReset) begin
      _T_1681 <= 4'h0;
    end else if (_T_1715) begin
      _T_1681 <= io_in_d_bits_size;
    end
    if (metaReset) begin
      _T_1683 <= 1'h0;
    end else if (_T_1715) begin
      _T_1683 <= io_in_d_bits_source;
    end
    if (metaReset) begin
      _T_1685 <= 2'h0;
    end else if (_T_1715) begin
      _T_1685 <= io_in_d_bits_sink;
    end
    if (metaReset) begin
      _T_1687 <= 1'h0;
    end else if (_T_1715) begin
      _T_1687 <= io_in_d_bits_denied;
    end
    if (metaReset) begin
      _T_1726 <= 9'h0;
    end else if (reset) begin
      _T_1726 <= 9'h0;
    end else if (_T_1716) begin
      if (_T_1730) begin
        _T_1726 <= 9'h0;
      end else begin
        _T_1726 <= _T_1729;
      end
    end
    if (metaReset) begin
      _T_1739 <= 3'h0;
    end else if (_T_1771) begin
      _T_1739 <= io_in_b_bits_opcode;
    end
    if (metaReset) begin
      _T_1741 <= 2'h0;
    end else if (_T_1771) begin
      _T_1741 <= io_in_b_bits_param;
    end
    if (metaReset) begin
      _T_1743 <= 4'h0;
    end else if (_T_1771) begin
      _T_1743 <= io_in_b_bits_size;
    end
    if (metaReset) begin
      _T_1745 <= 1'h0;
    end else if (_T_1771) begin
      _T_1745 <= io_in_b_bits_source;
    end
    if (metaReset) begin
      _T_1747 <= 32'h0;
    end else if (_T_1771) begin
      _T_1747 <= io_in_b_bits_address;
    end
    if (metaReset) begin
      _T_1781 <= 9'h0;
    end else if (reset) begin
      _T_1781 <= 9'h0;
    end else if (_T_1772) begin
      if (_T_1785) begin
        if (io_in_c_bits_opcode[0]) begin
          _T_1781 <= _T_1777;
        end else begin
          _T_1781 <= 9'h0;
        end
      end else begin
        _T_1781 <= _T_1784;
      end
    end
    if (metaReset) begin
      _T_1794 <= 3'h0;
    end else if (_T_1826) begin
      _T_1794 <= io_in_c_bits_opcode;
    end
    if (metaReset) begin
      _T_1796 <= 3'h0;
    end else if (_T_1826) begin
      _T_1796 <= io_in_c_bits_param;
    end
    if (metaReset) begin
      _T_1798 <= 4'h0;
    end else if (_T_1826) begin
      _T_1798 <= io_in_c_bits_size;
    end
    if (metaReset) begin
      _T_1800 <= 1'h0;
    end else if (_T_1826) begin
      _T_1800 <= io_in_c_bits_source;
    end
    if (metaReset) begin
      _T_1802 <= 32'h0;
    end else if (_T_1826) begin
      _T_1802 <= io_in_c_bits_address;
    end
    if (metaReset) begin
      _T_1828 <= 2'h0;
    end else if (reset) begin
      _T_1828 <= 2'h0;
    end else begin
      _T_1828 <= _T_1908;
    end
    if (metaReset) begin
      _T_1839 <= 9'h0;
    end else if (reset) begin
      _T_1839 <= 9'h0;
    end else if (_T_1599) begin
      if (_T_1843) begin
        if (~io_in_a_bits_opcode[2]) begin
          _T_1839 <= _T_1604;
        end else begin
          _T_1839 <= 9'h0;
        end
      end else begin
        _T_1839 <= _T_1842;
      end
    end
    if (metaReset) begin
      _T_1860 <= 9'h0;
    end else if (reset) begin
      _T_1860 <= 9'h0;
    end else if (_T_1655) begin
      if (_T_1864) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1860 <= _T_1660;
        end else begin
          _T_1860 <= 9'h0;
        end
      end else begin
        _T_1860 <= _T_1863;
      end
    end
    if (metaReset) begin
      _T_1926 <= 4'h0;
    end else if (reset) begin
      _T_1926 <= 4'h0;
    end else begin
      _T_1926 <= _T_1978;
    end
    if (metaReset) begin
      _T_1936 <= 9'h0;
    end else if (reset) begin
      _T_1936 <= 9'h0;
    end else if (_T_1655) begin
      if (_T_1940) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1936 <= _T_1660;
        end else begin
          _T_1936 <= 9'h0;
        end
      end else begin
        _T_1936 <= _T_1939;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_36 & ~_T_172) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at HellaCache.scala:220:21)\n    at Monitor.scala:49 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquireBlock type unsupported by manager\" + extra)\n"); // @[Monitor.scala 49:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_36 & ~_T_172) begin
          $fatal; // @[Monitor.scala 49:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_36 & ~_T_192) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at HellaCache.scala:220:21)\n    at Monitor.scala:50 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquireBlock from a client which does not support Probe\" + extra)\n"); // @[Monitor.scala 50:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_36 & ~_T_192) begin
          $fatal; // @[Monitor.scala 50:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_36 & ~_T_195) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:51 assert (source_ok, \"'A' channel AcquireBlock carries invalid source ID\" + extra)\n"); // @[Monitor.scala 51:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_36 & ~_T_195) begin
          $fatal; // @[Monitor.scala 51:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_36 & ~_T_199) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at HellaCache.scala:220:21)\n    at Monitor.scala:52 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquireBlock smaller than a beat\" + extra)\n"); // @[Monitor.scala 52:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_36 & ~_T_199) begin
          $fatal; // @[Monitor.scala 52:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_36 & ~_T_202) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at HellaCache.scala:220:21)\n    at Monitor.scala:53 assert (is_aligned, \"'A' channel AcquireBlock address not aligned to size\" + extra)\n"); // @[Monitor.scala 53:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_36 & ~_T_202) begin
          $fatal; // @[Monitor.scala 53:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_36 & ~_T_206) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:54 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquireBlock carries invalid grow param\" + extra)\n"); // @[Monitor.scala 54:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_36 & ~_T_206) begin
          $fatal; // @[Monitor.scala 54:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_36 & ~_T_211) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at HellaCache.scala:220:21)\n    at Monitor.scala:55 assert (~bundle.mask === UInt(0), \"'A' channel AcquireBlock contains invalid mask\" + extra)\n"); // @[Monitor.scala 55:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_36 & ~_T_211) begin
          $fatal; // @[Monitor.scala 55:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_50 & ~_T_172) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at HellaCache.scala:220:21)\n    at Monitor.scala:60 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquirePerm type unsupported by manager\" + extra)\n"); // @[Monitor.scala 60:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_50 & ~_T_172) begin
          $fatal; // @[Monitor.scala 60:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_50 & ~_T_192) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at HellaCache.scala:220:21)\n    at Monitor.scala:61 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquirePerm from a client which does not support Probe\" + extra)\n"); // @[Monitor.scala 61:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_50 & ~_T_192) begin
          $fatal; // @[Monitor.scala 61:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_50 & ~_T_195) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:62 assert (source_ok, \"'A' channel AcquirePerm carries invalid source ID\" + extra)\n"); // @[Monitor.scala 62:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_50 & ~_T_195) begin
          $fatal; // @[Monitor.scala 62:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_50 & ~_T_199) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at HellaCache.scala:220:21)\n    at Monitor.scala:63 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquirePerm smaller than a beat\" + extra)\n"); // @[Monitor.scala 63:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_50 & ~_T_199) begin
          $fatal; // @[Monitor.scala 63:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_50 & ~_T_202) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at HellaCache.scala:220:21)\n    at Monitor.scala:64 assert (is_aligned, \"'A' channel AcquirePerm address not aligned to size\" + extra)\n"); // @[Monitor.scala 64:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_50 & ~_T_202) begin
          $fatal; // @[Monitor.scala 64:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_50 & ~_T_206) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:65 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquirePerm carries invalid grow param\" + extra)\n"); // @[Monitor.scala 65:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_50 & ~_T_206) begin
          $fatal; // @[Monitor.scala 65:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_50 & ~_T_306) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at HellaCache.scala:220:21)\n    at Monitor.scala:66 assert (bundle.param =/= TLPermissions.NtoB, \"'A' channel AcquirePerm requests NtoB\" + extra)\n"); // @[Monitor.scala 66:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_50 & ~_T_306) begin
          $fatal; // @[Monitor.scala 66:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_50 & ~_T_211) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at HellaCache.scala:220:21)\n    at Monitor.scala:67 assert (~bundle.mask === UInt(0), \"'A' channel AcquirePerm contains invalid mask\" + extra)\n"); // @[Monitor.scala 67:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_50 & ~_T_211) begin
          $fatal; // @[Monitor.scala 67:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_66 & ~_T_371) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at HellaCache.scala:220:21)\n    at Monitor.scala:72 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); // @[Monitor.scala 72:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_66 & ~_T_371) begin
          $fatal; // @[Monitor.scala 72:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_66 & ~_T_195) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:73 assert (source_ok, \"'A' channel Get carries invalid source ID\" + extra)\n"); // @[Monitor.scala 73:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_66 & ~_T_195) begin
          $fatal; // @[Monitor.scala 73:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_66 & ~_T_202) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at HellaCache.scala:220:21)\n    at Monitor.scala:74 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); // @[Monitor.scala 74:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_66 & ~_T_202) begin
          $fatal; // @[Monitor.scala 74:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_66 & ~_T_381) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:75 assert (bundle.param === UInt(0), \"'A' channel Get carries invalid param\" + extra)\n"); // @[Monitor.scala 75:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_66 & ~_T_381) begin
          $fatal; // @[Monitor.scala 75:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_66 & ~_T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at HellaCache.scala:220:21)\n    at Monitor.scala:76 assert (bundle.mask === mask, \"'A' channel Get contains invalid mask\" + extra)\n"); // @[Monitor.scala 76:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_66 & ~_T_385) begin
          $fatal; // @[Monitor.scala 76:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_76 & ~_T_452) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at HellaCache.scala:220:21)\n    at Monitor.scala:81 assert (edge.manager.supportsPutFullSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutFull type unsupported by manager\" + extra)\n"); // @[Monitor.scala 81:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_76 & ~_T_452) begin
          $fatal; // @[Monitor.scala 81:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_76 & ~_T_195) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:82 assert (source_ok, \"'A' channel PutFull carries invalid source ID\" + extra)\n"); // @[Monitor.scala 82:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_76 & ~_T_195) begin
          $fatal; // @[Monitor.scala 82:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_76 & ~_T_202) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at HellaCache.scala:220:21)\n    at Monitor.scala:83 assert (is_aligned, \"'A' channel PutFull address not aligned to size\" + extra)\n"); // @[Monitor.scala 83:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_76 & ~_T_202) begin
          $fatal; // @[Monitor.scala 83:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_76 & ~_T_381) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:84 assert (bundle.param === UInt(0), \"'A' channel PutFull carries invalid param\" + extra)\n"); // @[Monitor.scala 84:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_76 & ~_T_381) begin
          $fatal; // @[Monitor.scala 84:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_76 & ~_T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at HellaCache.scala:220:21)\n    at Monitor.scala:85 assert (bundle.mask === mask, \"'A' channel PutFull contains invalid mask\" + extra)\n"); // @[Monitor.scala 85:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_76 & ~_T_385) begin
          $fatal; // @[Monitor.scala 85:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_86 & ~_T_452) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at HellaCache.scala:220:21)\n    at Monitor.scala:89 assert (edge.manager.supportsPutPartialSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutPartial type unsupported by manager\" + extra)\n"); // @[Monitor.scala 89:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_86 & ~_T_452) begin
          $fatal; // @[Monitor.scala 89:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_86 & ~_T_195) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:90 assert (source_ok, \"'A' channel PutPartial carries invalid source ID\" + extra)\n"); // @[Monitor.scala 90:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_86 & ~_T_195) begin
          $fatal; // @[Monitor.scala 90:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_86 & ~_T_202) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at HellaCache.scala:220:21)\n    at Monitor.scala:91 assert (is_aligned, \"'A' channel PutPartial address not aligned to size\" + extra)\n"); // @[Monitor.scala 91:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_86 & ~_T_202) begin
          $fatal; // @[Monitor.scala 91:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_86 & ~_T_381) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:92 assert (bundle.param === UInt(0), \"'A' channel PutPartial carries invalid param\" + extra)\n"); // @[Monitor.scala 92:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_86 & ~_T_381) begin
          $fatal; // @[Monitor.scala 92:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_86 & ~_T_545) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at HellaCache.scala:220:21)\n    at Monitor.scala:93 assert ((bundle.mask & ~mask) === UInt(0), \"'A' channel PutPartial contains invalid mask\" + extra)\n"); // @[Monitor.scala 93:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_86 & ~_T_545) begin
          $fatal; // @[Monitor.scala 93:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_96 & ~_T_598) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at HellaCache.scala:220:21)\n    at Monitor.scala:97 assert (edge.manager.supportsArithmeticSafe(edge.address(bundle), bundle.size), \"'A' channel carries Arithmetic type unsupported by manager\" + extra)\n"); // @[Monitor.scala 97:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_96 & ~_T_598) begin
          $fatal; // @[Monitor.scala 97:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_96 & ~_T_195) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:98 assert (source_ok, \"'A' channel Arithmetic carries invalid source ID\" + extra)\n"); // @[Monitor.scala 98:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_96 & ~_T_195) begin
          $fatal; // @[Monitor.scala 98:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_96 & ~_T_202) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at HellaCache.scala:220:21)\n    at Monitor.scala:99 assert (is_aligned, \"'A' channel Arithmetic address not aligned to size\" + extra)\n"); // @[Monitor.scala 99:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_96 & ~_T_202) begin
          $fatal; // @[Monitor.scala 99:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_96 & ~_T_608) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:100 assert (TLAtomics.isArithmetic(bundle.param), \"'A' channel Arithmetic carries invalid opcode param\" + extra)\n"); // @[Monitor.scala 100:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_96 & ~_T_608) begin
          $fatal; // @[Monitor.scala 100:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_96 & ~_T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at HellaCache.scala:220:21)\n    at Monitor.scala:101 assert (bundle.mask === mask, \"'A' channel Arithmetic contains invalid mask\" + extra)\n"); // @[Monitor.scala 101:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_96 & ~_T_385) begin
          $fatal; // @[Monitor.scala 101:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_106 & ~_T_598) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at HellaCache.scala:220:21)\n    at Monitor.scala:105 assert (edge.manager.supportsLogicalSafe(edge.address(bundle), bundle.size), \"'A' channel carries Logical type unsupported by manager\" + extra)\n"); // @[Monitor.scala 105:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_106 & ~_T_598) begin
          $fatal; // @[Monitor.scala 105:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_106 & ~_T_195) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:106 assert (source_ok, \"'A' channel Logical carries invalid source ID\" + extra)\n"); // @[Monitor.scala 106:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_106 & ~_T_195) begin
          $fatal; // @[Monitor.scala 106:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_106 & ~_T_202) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at HellaCache.scala:220:21)\n    at Monitor.scala:107 assert (is_aligned, \"'A' channel Logical address not aligned to size\" + extra)\n"); // @[Monitor.scala 107:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_106 & ~_T_202) begin
          $fatal; // @[Monitor.scala 107:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_106 & ~_T_675) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:108 assert (TLAtomics.isLogical(bundle.param), \"'A' channel Logical carries invalid opcode param\" + extra)\n"); // @[Monitor.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_106 & ~_T_675) begin
          $fatal; // @[Monitor.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_106 & ~_T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at HellaCache.scala:220:21)\n    at Monitor.scala:109 assert (bundle.mask === mask, \"'A' channel Logical contains invalid mask\" + extra)\n"); // @[Monitor.scala 109:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_106 & ~_T_385) begin
          $fatal; // @[Monitor.scala 109:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_116 & ~_T_732) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at HellaCache.scala:220:21)\n    at Monitor.scala:113 assert (edge.manager.supportsHintSafe(edge.address(bundle), bundle.size), \"'A' channel carries Hint type unsupported by manager\" + extra)\n"); // @[Monitor.scala 113:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_116 & ~_T_732) begin
          $fatal; // @[Monitor.scala 113:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_116 & ~_T_195) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:114 assert (source_ok, \"'A' channel Hint carries invalid source ID\" + extra)\n"); // @[Monitor.scala 114:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_116 & ~_T_195) begin
          $fatal; // @[Monitor.scala 114:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_116 & ~_T_202) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at HellaCache.scala:220:21)\n    at Monitor.scala:115 assert (is_aligned, \"'A' channel Hint address not aligned to size\" + extra)\n"); // @[Monitor.scala 115:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_116 & ~_T_202) begin
          $fatal; // @[Monitor.scala 115:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_116 & ~_T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at HellaCache.scala:220:21)\n    at Monitor.scala:116 assert (bundle.mask === mask, \"'A' channel Hint contains invalid mask\" + extra)\n"); // @[Monitor.scala 116:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_116 & ~_T_385) begin
          $fatal; // @[Monitor.scala 116:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~_T_750) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at HellaCache.scala:220:21)\n    at Monitor.scala:268 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); // @[Monitor.scala 268:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~_T_750) begin
          $fatal; // @[Monitor.scala 268:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_124 & ~_T_766) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:276 assert (source_ok, \"'D' channel ReleaseAck carries invalid source ID\" + extra)\n"); // @[Monitor.scala 276:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_124 & ~_T_766) begin
          $fatal; // @[Monitor.scala 276:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_124 & ~_T_770) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at HellaCache.scala:220:21)\n    at Monitor.scala:277 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); // @[Monitor.scala 277:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_124 & ~_T_770) begin
          $fatal; // @[Monitor.scala 277:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_124 & ~_T_774) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:278 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); // @[Monitor.scala 278:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_124 & ~_T_774) begin
          $fatal; // @[Monitor.scala 278:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_124 & ~_T_778) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at HellaCache.scala:220:21)\n    at Monitor.scala:279 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); // @[Monitor.scala 279:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_124 & ~_T_778) begin
          $fatal; // @[Monitor.scala 279:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_124 & ~_T_782) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at HellaCache.scala:220:21)\n    at Monitor.scala:280 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); // @[Monitor.scala 280:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_124 & ~_T_782) begin
          $fatal; // @[Monitor.scala 280:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_134 & ~_T_766) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:284 assert (source_ok, \"'D' channel Grant carries invalid source ID\" + extra)\n"); // @[Monitor.scala 284:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_134 & ~_T_766) begin
          $fatal; // @[Monitor.scala 284:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_134 & ~_T_770) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at HellaCache.scala:220:21)\n    at Monitor.scala:286 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); // @[Monitor.scala 286:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_134 & ~_T_770) begin
          $fatal; // @[Monitor.scala 286:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_134 & ~_T_797) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:287 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); // @[Monitor.scala 287:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_134 & ~_T_797) begin
          $fatal; // @[Monitor.scala 287:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_134 & ~_T_801) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:288 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); // @[Monitor.scala 288:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_134 & ~_T_801) begin
          $fatal; // @[Monitor.scala 288:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_134 & ~_T_778) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at HellaCache.scala:220:21)\n    at Monitor.scala:289 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); // @[Monitor.scala 289:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_134 & ~_T_778) begin
          $fatal; // @[Monitor.scala 289:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & ~_T_766) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:294 assert (source_ok, \"'D' channel GrantData carries invalid source ID\" + extra)\n"); // @[Monitor.scala 294:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & ~_T_766) begin
          $fatal; // @[Monitor.scala 294:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & ~_T_770) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at HellaCache.scala:220:21)\n    at Monitor.scala:296 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); // @[Monitor.scala 296:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & ~_T_770) begin
          $fatal; // @[Monitor.scala 296:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & ~_T_797) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:297 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); // @[Monitor.scala 297:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & ~_T_797) begin
          $fatal; // @[Monitor.scala 297:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & ~_T_801) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:298 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); // @[Monitor.scala 298:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & ~_T_801) begin
          $fatal; // @[Monitor.scala 298:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & ~_T_834) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at HellaCache.scala:220:21)\n    at Monitor.scala:299 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); // @[Monitor.scala 299:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & ~_T_834) begin
          $fatal; // @[Monitor.scala 299:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_154 & ~_T_766) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:304 assert (source_ok, \"'D' channel AccessAck carries invalid source ID\" + extra)\n"); // @[Monitor.scala 304:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_154 & ~_T_766) begin
          $fatal; // @[Monitor.scala 304:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_154 & ~_T_774) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:306 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); // @[Monitor.scala 306:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_154 & ~_T_774) begin
          $fatal; // @[Monitor.scala 306:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_154 & ~_T_778) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at HellaCache.scala:220:21)\n    at Monitor.scala:307 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); // @[Monitor.scala 307:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_154 & ~_T_778) begin
          $fatal; // @[Monitor.scala 307:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & ~_T_766) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:312 assert (source_ok, \"'D' channel AccessAckData carries invalid source ID\" + extra)\n"); // @[Monitor.scala 312:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & ~_T_766) begin
          $fatal; // @[Monitor.scala 312:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & ~_T_774) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:314 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); // @[Monitor.scala 314:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & ~_T_774) begin
          $fatal; // @[Monitor.scala 314:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & ~_T_834) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at HellaCache.scala:220:21)\n    at Monitor.scala:315 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); // @[Monitor.scala 315:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & ~_T_834) begin
          $fatal; // @[Monitor.scala 315:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & ~_T_766) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:320 assert (source_ok, \"'D' channel HintAck carries invalid source ID\" + extra)\n"); // @[Monitor.scala 320:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & ~_T_766) begin
          $fatal; // @[Monitor.scala 320:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & ~_T_774) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:322 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); // @[Monitor.scala 322:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & ~_T_774) begin
          $fatal; // @[Monitor.scala 322:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & ~_T_778) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at HellaCache.scala:220:21)\n    at Monitor.scala:323 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); // @[Monitor.scala 323:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & ~_T_778) begin
          $fatal; // @[Monitor.scala 323:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_b_valid & ~_T_895) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel has invalid opcode (connected at HellaCache.scala:220:21)\n    at Monitor.scala:122 assert (TLMessages.isB(bundle.opcode), \"'B' channel has invalid opcode\" + extra)\n"); // @[Monitor.scala 122:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_b_valid & ~_T_895) begin
          $fatal; // @[Monitor.scala 122:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_172 & ~_T_1077) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Probe type unsupported by client (connected at HellaCache.scala:220:21)\n    at Monitor.scala:133 assert (edge.client.supportsProbe(bundle.source, bundle.size), \"'B' channel carries Probe type unsupported by client\" + extra)\n"); // @[Monitor.scala 133:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_172 & ~_T_1077) begin
          $fatal; // @[Monitor.scala 133:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_172 & ~_T_1080) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries unmanaged address (connected at HellaCache.scala:220:21)\n    at Monitor.scala:134 assert (address_ok, \"'B' channel Probe carries unmanaged address\" + extra)\n"); // @[Monitor.scala 134:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_172 & ~_T_1080) begin
          $fatal; // @[Monitor.scala 134:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_172 & ~_T_1083) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries source that is not first source (connected at HellaCache.scala:220:21)\n    at Monitor.scala:135 assert (legal_source, \"'B' channel Probe carries source that is not first source\" + extra)\n"); // @[Monitor.scala 135:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_172 & ~_T_1083) begin
          $fatal; // @[Monitor.scala 135:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_172 & ~_T_1086) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe address not aligned to size (connected at HellaCache.scala:220:21)\n    at Monitor.scala:136 assert (is_aligned, \"'B' channel Probe address not aligned to size\" + extra)\n"); // @[Monitor.scala 136:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_172 & ~_T_1086) begin
          $fatal; // @[Monitor.scala 136:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_172 & ~_T_1090) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries invalid cap param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:137 assert (TLPermissions.isCap(bundle.param), \"'B' channel Probe carries invalid cap param\" + extra)\n"); // @[Monitor.scala 137:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_172 & ~_T_1090) begin
          $fatal; // @[Monitor.scala 137:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_172 & ~_T_1094) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe contains invalid mask (connected at HellaCache.scala:220:21)\n    at Monitor.scala:138 assert (bundle.mask === mask, \"'B' channel Probe contains invalid mask\" + extra)\n"); // @[Monitor.scala 138:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_172 & ~_T_1094) begin
          $fatal; // @[Monitor.scala 138:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_172 & ~_T_1098) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe is corrupt (connected at HellaCache.scala:220:21)\n    at Monitor.scala:139 assert (!bundle.corrupt, \"'B' channel Probe is corrupt\" + extra)\n"); // @[Monitor.scala 139:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_172 & ~_T_1098) begin
          $fatal; // @[Monitor.scala 139:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Get type unsupported by client (connected at HellaCache.scala:220:21)\n    at Monitor.scala:143 assert (edge.client.supportsGet(bundle.source, bundle.size), \"'B' channel carries Get type unsupported by client\" + extra)\n"); // @[Monitor.scala 143:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & ~reset) begin
          $fatal; // @[Monitor.scala 143:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & ~_T_1080) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries unmanaged address (connected at HellaCache.scala:220:21)\n    at Monitor.scala:144 assert (address_ok, \"'B' channel Get carries unmanaged address\" + extra)\n"); // @[Monitor.scala 144:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & ~_T_1080) begin
          $fatal; // @[Monitor.scala 144:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & ~_T_1083) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries source that is not first source (connected at HellaCache.scala:220:21)\n    at Monitor.scala:145 assert (legal_source, \"'B' channel Get carries source that is not first source\" + extra)\n"); // @[Monitor.scala 145:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & ~_T_1083) begin
          $fatal; // @[Monitor.scala 145:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & ~_T_1086) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get address not aligned to size (connected at HellaCache.scala:220:21)\n    at Monitor.scala:146 assert (is_aligned, \"'B' channel Get address not aligned to size\" + extra)\n"); // @[Monitor.scala 146:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & ~_T_1086) begin
          $fatal; // @[Monitor.scala 146:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & ~_T_1115) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries invalid param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:147 assert (bundle.param === UInt(0), \"'B' channel Get carries invalid param\" + extra)\n"); // @[Monitor.scala 147:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & ~_T_1115) begin
          $fatal; // @[Monitor.scala 147:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & ~_T_1094) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get contains invalid mask (connected at HellaCache.scala:220:21)\n    at Monitor.scala:148 assert (bundle.mask === mask, \"'B' channel Get contains invalid mask\" + extra)\n"); // @[Monitor.scala 148:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & ~_T_1094) begin
          $fatal; // @[Monitor.scala 148:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & ~_T_1098) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get is corrupt (connected at HellaCache.scala:220:21)\n    at Monitor.scala:149 assert (!bundle.corrupt, \"'B' channel Get is corrupt\" + extra)\n"); // @[Monitor.scala 149:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & ~_T_1098) begin
          $fatal; // @[Monitor.scala 149:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_200 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutFull type unsupported by client (connected at HellaCache.scala:220:21)\n    at Monitor.scala:153 assert (edge.client.supportsPutFull(bundle.source, bundle.size), \"'B' channel carries PutFull type unsupported by client\" + extra)\n"); // @[Monitor.scala 153:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_200 & ~reset) begin
          $fatal; // @[Monitor.scala 153:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_200 & ~_T_1080) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries unmanaged address (connected at HellaCache.scala:220:21)\n    at Monitor.scala:154 assert (address_ok, \"'B' channel PutFull carries unmanaged address\" + extra)\n"); // @[Monitor.scala 154:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_200 & ~_T_1080) begin
          $fatal; // @[Monitor.scala 154:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_200 & ~_T_1083) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries source that is not first source (connected at HellaCache.scala:220:21)\n    at Monitor.scala:155 assert (legal_source, \"'B' channel PutFull carries source that is not first source\" + extra)\n"); // @[Monitor.scala 155:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_200 & ~_T_1083) begin
          $fatal; // @[Monitor.scala 155:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_200 & ~_T_1086) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull address not aligned to size (connected at HellaCache.scala:220:21)\n    at Monitor.scala:156 assert (is_aligned, \"'B' channel PutFull address not aligned to size\" + extra)\n"); // @[Monitor.scala 156:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_200 & ~_T_1086) begin
          $fatal; // @[Monitor.scala 156:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_200 & ~_T_1115) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries invalid param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:157 assert (bundle.param === UInt(0), \"'B' channel PutFull carries invalid param\" + extra)\n"); // @[Monitor.scala 157:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_200 & ~_T_1115) begin
          $fatal; // @[Monitor.scala 157:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_200 & ~_T_1094) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull contains invalid mask (connected at HellaCache.scala:220:21)\n    at Monitor.scala:158 assert (bundle.mask === mask, \"'B' channel PutFull contains invalid mask\" + extra)\n"); // @[Monitor.scala 158:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_200 & ~_T_1094) begin
          $fatal; // @[Monitor.scala 158:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_212 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutPartial type unsupported by client (connected at HellaCache.scala:220:21)\n    at Monitor.scala:162 assert (edge.client.supportsPutPartial(bundle.source, bundle.size), \"'B' channel carries PutPartial type unsupported by client\" + extra)\n"); // @[Monitor.scala 162:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_212 & ~reset) begin
          $fatal; // @[Monitor.scala 162:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_212 & ~_T_1080) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at HellaCache.scala:220:21)\n    at Monitor.scala:163 assert (address_ok, \"'B' channel PutPartial carries unmanaged address\" + extra)\n"); // @[Monitor.scala 163:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_212 & ~_T_1080) begin
          $fatal; // @[Monitor.scala 163:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_212 & ~_T_1083) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries source that is not first source (connected at HellaCache.scala:220:21)\n    at Monitor.scala:164 assert (legal_source, \"'B' channel PutPartial carries source that is not first source\" + extra)\n"); // @[Monitor.scala 164:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_212 & ~_T_1083) begin
          $fatal; // @[Monitor.scala 164:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_212 & ~_T_1086) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial address not aligned to size (connected at HellaCache.scala:220:21)\n    at Monitor.scala:165 assert (is_aligned, \"'B' channel PutPartial address not aligned to size\" + extra)\n"); // @[Monitor.scala 165:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_212 & ~_T_1086) begin
          $fatal; // @[Monitor.scala 165:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_212 & ~_T_1115) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries invalid param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:166 assert (bundle.param === UInt(0), \"'B' channel PutPartial carries invalid param\" + extra)\n"); // @[Monitor.scala 166:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_212 & ~_T_1115) begin
          $fatal; // @[Monitor.scala 166:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_212 & ~_T_1167) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial contains invalid mask (connected at HellaCache.scala:220:21)\n    at Monitor.scala:167 assert ((bundle.mask & ~mask) === UInt(0), \"'B' channel PutPartial contains invalid mask\" + extra)\n"); // @[Monitor.scala 167:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_212 & ~_T_1167) begin
          $fatal; // @[Monitor.scala 167:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_224 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Arithmetic type unsupported by client (connected at HellaCache.scala:220:21)\n    at Monitor.scala:171 assert (edge.client.supportsArithmetic(bundle.source, bundle.size), \"'B' channel carries Arithmetic type unsupported by client\" + extra)\n"); // @[Monitor.scala 171:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_224 & ~reset) begin
          $fatal; // @[Monitor.scala 171:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_224 & ~_T_1080) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at HellaCache.scala:220:21)\n    at Monitor.scala:172 assert (address_ok, \"'B' channel Arithmetic carries unmanaged address\" + extra)\n"); // @[Monitor.scala 172:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_224 & ~_T_1080) begin
          $fatal; // @[Monitor.scala 172:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_224 & ~_T_1083) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries source that is not first source (connected at HellaCache.scala:220:21)\n    at Monitor.scala:173 assert (legal_source, \"'B' channel Arithmetic carries source that is not first source\" + extra)\n"); // @[Monitor.scala 173:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_224 & ~_T_1083) begin
          $fatal; // @[Monitor.scala 173:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_224 & ~_T_1086) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at HellaCache.scala:220:21)\n    at Monitor.scala:174 assert (is_aligned, \"'B' channel Arithmetic address not aligned to size\" + extra)\n"); // @[Monitor.scala 174:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_224 & ~_T_1086) begin
          $fatal; // @[Monitor.scala 174:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_224 & ~_T_1094) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at HellaCache.scala:220:21)\n    at Monitor.scala:176 assert (bundle.mask === mask, \"'B' channel Arithmetic contains invalid mask\" + extra)\n"); // @[Monitor.scala 176:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_224 & ~_T_1094) begin
          $fatal; // @[Monitor.scala 176:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_234 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Logical type unsupported by client (connected at HellaCache.scala:220:21)\n    at Monitor.scala:180 assert (edge.client.supportsLogical(bundle.source, bundle.size), \"'B' channel carries Logical type unsupported by client\" + extra)\n"); // @[Monitor.scala 180:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_234 & ~reset) begin
          $fatal; // @[Monitor.scala 180:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_234 & ~_T_1080) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries unmanaged address (connected at HellaCache.scala:220:21)\n    at Monitor.scala:181 assert (address_ok, \"'B' channel Logical carries unmanaged address\" + extra)\n"); // @[Monitor.scala 181:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_234 & ~_T_1080) begin
          $fatal; // @[Monitor.scala 181:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_234 & ~_T_1083) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries source that is not first source (connected at HellaCache.scala:220:21)\n    at Monitor.scala:182 assert (legal_source, \"'B' channel Logical carries source that is not first source\" + extra)\n"); // @[Monitor.scala 182:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_234 & ~_T_1083) begin
          $fatal; // @[Monitor.scala 182:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_234 & ~_T_1086) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical address not aligned to size (connected at HellaCache.scala:220:21)\n    at Monitor.scala:183 assert (is_aligned, \"'B' channel Logical address not aligned to size\" + extra)\n"); // @[Monitor.scala 183:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_234 & ~_T_1086) begin
          $fatal; // @[Monitor.scala 183:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_234 & ~_T_1094) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical contains invalid mask (connected at HellaCache.scala:220:21)\n    at Monitor.scala:185 assert (bundle.mask === mask, \"'B' channel Logical contains invalid mask\" + extra)\n"); // @[Monitor.scala 185:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_234 & ~_T_1094) begin
          $fatal; // @[Monitor.scala 185:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Hint type unsupported by client (connected at HellaCache.scala:220:21)\n    at Monitor.scala:189 assert (edge.client.supportsHint(bundle.source, bundle.size), \"'B' channel carries Hint type unsupported by client\" + extra)\n"); // @[Monitor.scala 189:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & ~reset) begin
          $fatal; // @[Monitor.scala 189:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & ~_T_1080) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries unmanaged address (connected at HellaCache.scala:220:21)\n    at Monitor.scala:190 assert (address_ok, \"'B' channel Hint carries unmanaged address\" + extra)\n"); // @[Monitor.scala 190:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & ~_T_1080) begin
          $fatal; // @[Monitor.scala 190:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & ~_T_1083) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries source that is not first source (connected at HellaCache.scala:220:21)\n    at Monitor.scala:191 assert (legal_source, \"'B' channel Hint carries source that is not first source\" + extra)\n"); // @[Monitor.scala 191:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & ~_T_1083) begin
          $fatal; // @[Monitor.scala 191:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & ~_T_1086) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint address not aligned to size (connected at HellaCache.scala:220:21)\n    at Monitor.scala:192 assert (is_aligned, \"'B' channel Hint address not aligned to size\" + extra)\n"); // @[Monitor.scala 192:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & ~_T_1086) begin
          $fatal; // @[Monitor.scala 192:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & ~_T_1094) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint contains invalid mask (connected at HellaCache.scala:220:21)\n    at Monitor.scala:193 assert (bundle.mask === mask, \"'B' channel Hint contains invalid mask\" + extra)\n"); // @[Monitor.scala 193:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & ~_T_1094) begin
          $fatal; // @[Monitor.scala 193:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & ~_T_1098) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint is corrupt (connected at HellaCache.scala:220:21)\n    at Monitor.scala:194 assert (!bundle.corrupt, \"'B' channel Hint is corrupt\" + extra)\n"); // @[Monitor.scala 194:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & ~_T_1098) begin
          $fatal; // @[Monitor.scala 194:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_256 & ~_T_1329) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at HellaCache.scala:220:21)\n    at Monitor.scala:208 assert (address_ok, \"'C' channel ProbeAck carries unmanaged address\" + extra)\n"); // @[Monitor.scala 208:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_256 & ~_T_1329) begin
          $fatal; // @[Monitor.scala 208:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_256 & ~_T_1332) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:209 assert (source_ok, \"'C' channel ProbeAck carries invalid source ID\" + extra)\n"); // @[Monitor.scala 209:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_256 & ~_T_1332) begin
          $fatal; // @[Monitor.scala 209:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_256 & ~_T_1336) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at HellaCache.scala:220:21)\n    at Monitor.scala:210 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAck smaller than a beat\" + extra)\n"); // @[Monitor.scala 210:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_256 & ~_T_1336) begin
          $fatal; // @[Monitor.scala 210:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_256 & ~_T_1339) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at HellaCache.scala:220:21)\n    at Monitor.scala:211 assert (is_aligned, \"'C' channel ProbeAck address not aligned to size\" + extra)\n"); // @[Monitor.scala 211:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_256 & ~_T_1339) begin
          $fatal; // @[Monitor.scala 211:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_256 & ~_T_1343) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:212 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAck carries invalid report param\" + extra)\n"); // @[Monitor.scala 212:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_256 & ~_T_1343) begin
          $fatal; // @[Monitor.scala 212:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_266 & ~_T_1329) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at HellaCache.scala:220:21)\n    at Monitor.scala:217 assert (address_ok, \"'C' channel ProbeAckData carries unmanaged address\" + extra)\n"); // @[Monitor.scala 217:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_266 & ~_T_1329) begin
          $fatal; // @[Monitor.scala 217:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_266 & ~_T_1332) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:218 assert (source_ok, \"'C' channel ProbeAckData carries invalid source ID\" + extra)\n"); // @[Monitor.scala 218:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_266 & ~_T_1332) begin
          $fatal; // @[Monitor.scala 218:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_266 & ~_T_1336) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at HellaCache.scala:220:21)\n    at Monitor.scala:219 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAckData smaller than a beat\" + extra)\n"); // @[Monitor.scala 219:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_266 & ~_T_1336) begin
          $fatal; // @[Monitor.scala 219:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_266 & ~_T_1339) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at HellaCache.scala:220:21)\n    at Monitor.scala:220 assert (is_aligned, \"'C' channel ProbeAckData address not aligned to size\" + extra)\n"); // @[Monitor.scala 220:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_266 & ~_T_1339) begin
          $fatal; // @[Monitor.scala 220:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_266 & ~_T_1343) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:221 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAckData carries invalid report param\" + extra)\n"); // @[Monitor.scala 221:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_266 & ~_T_1343) begin
          $fatal; // @[Monitor.scala 221:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_276 & ~_T_1418) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release type unsupported by manager (connected at HellaCache.scala:220:21)\n    at Monitor.scala:225 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries Release type unsupported by manager\" + extra)\n"); // @[Monitor.scala 225:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_276 & ~_T_1418) begin
          $fatal; // @[Monitor.scala 225:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_276 & ~_T_1438) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at HellaCache.scala:220:21)\n    at Monitor.scala:226 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); // @[Monitor.scala 226:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_276 & ~_T_1438) begin
          $fatal; // @[Monitor.scala 226:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_276 & ~_T_1332) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid source ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:227 assert (source_ok, \"'C' channel Release carries invalid source ID\" + extra)\n"); // @[Monitor.scala 227:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_276 & ~_T_1332) begin
          $fatal; // @[Monitor.scala 227:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_276 & ~_T_1336) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release smaller than a beat (connected at HellaCache.scala:220:21)\n    at Monitor.scala:228 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel Release smaller than a beat\" + extra)\n"); // @[Monitor.scala 228:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_276 & ~_T_1336) begin
          $fatal; // @[Monitor.scala 228:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_276 & ~_T_1339) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release address not aligned to size (connected at HellaCache.scala:220:21)\n    at Monitor.scala:229 assert (is_aligned, \"'C' channel Release address not aligned to size\" + extra)\n"); // @[Monitor.scala 229:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_276 & ~_T_1339) begin
          $fatal; // @[Monitor.scala 229:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_276 & ~_T_1452) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid shrink param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:230 assert (TLPermissions.isShrink(bundle.param), \"'C' channel Release carries invalid shrink param\" + extra)\n"); // @[Monitor.scala 230:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_276 & ~_T_1452) begin
          $fatal; // @[Monitor.scala 230:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_288 & ~_T_1418) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at HellaCache.scala:220:21)\n    at Monitor.scala:235 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries ReleaseData type unsupported by manager\" + extra)\n"); // @[Monitor.scala 235:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_288 & ~_T_1418) begin
          $fatal; // @[Monitor.scala 235:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_288 & ~_T_1438) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at HellaCache.scala:220:21)\n    at Monitor.scala:236 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); // @[Monitor.scala 236:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_288 & ~_T_1438) begin
          $fatal; // @[Monitor.scala 236:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_288 & ~_T_1332) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:237 assert (source_ok, \"'C' channel ReleaseData carries invalid source ID\" + extra)\n"); // @[Monitor.scala 237:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_288 & ~_T_1332) begin
          $fatal; // @[Monitor.scala 237:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_288 & ~_T_1336) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at HellaCache.scala:220:21)\n    at Monitor.scala:238 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ReleaseData smaller than a beat\" + extra)\n"); // @[Monitor.scala 238:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_288 & ~_T_1336) begin
          $fatal; // @[Monitor.scala 238:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_288 & ~_T_1339) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at HellaCache.scala:220:21)\n    at Monitor.scala:239 assert (is_aligned, \"'C' channel ReleaseData address not aligned to size\" + extra)\n"); // @[Monitor.scala 239:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_288 & ~_T_1339) begin
          $fatal; // @[Monitor.scala 239:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_288 & ~_T_1452) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid shrink param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:240 assert (TLPermissions.isShrink(bundle.param), \"'C' channel ReleaseData carries invalid shrink param\" + extra)\n"); // @[Monitor.scala 240:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_288 & ~_T_1452) begin
          $fatal; // @[Monitor.scala 240:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_300 & ~_T_1329) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at HellaCache.scala:220:21)\n    at Monitor.scala:244 assert (address_ok, \"'C' channel AccessAck carries unmanaged address\" + extra)\n"); // @[Monitor.scala 244:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_300 & ~_T_1329) begin
          $fatal; // @[Monitor.scala 244:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_300 & ~_T_1332) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:245 assert (source_ok, \"'C' channel AccessAck carries invalid source ID\" + extra)\n"); // @[Monitor.scala 245:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_300 & ~_T_1332) begin
          $fatal; // @[Monitor.scala 245:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_300 & ~_T_1339) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck address not aligned to size (connected at HellaCache.scala:220:21)\n    at Monitor.scala:246 assert (is_aligned, \"'C' channel AccessAck address not aligned to size\" + extra)\n"); // @[Monitor.scala 246:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_300 & ~_T_1339) begin
          $fatal; // @[Monitor.scala 246:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_300 & ~_T_1557) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:247 assert (bundle.param === UInt(0), \"'C' channel AccessAck carries invalid param\" + extra)\n"); // @[Monitor.scala 247:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_300 & ~_T_1557) begin
          $fatal; // @[Monitor.scala 247:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_308 & ~_T_1329) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at HellaCache.scala:220:21)\n    at Monitor.scala:252 assert (address_ok, \"'C' channel AccessAckData carries unmanaged address\" + extra)\n"); // @[Monitor.scala 252:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_308 & ~_T_1329) begin
          $fatal; // @[Monitor.scala 252:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_308 & ~_T_1332) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:253 assert (source_ok, \"'C' channel AccessAckData carries invalid source ID\" + extra)\n"); // @[Monitor.scala 253:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_308 & ~_T_1332) begin
          $fatal; // @[Monitor.scala 253:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_308 & ~_T_1339) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at HellaCache.scala:220:21)\n    at Monitor.scala:254 assert (is_aligned, \"'C' channel AccessAckData address not aligned to size\" + extra)\n"); // @[Monitor.scala 254:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_308 & ~_T_1339) begin
          $fatal; // @[Monitor.scala 254:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_308 & ~_T_1557) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:255 assert (bundle.param === UInt(0), \"'C' channel AccessAckData carries invalid param\" + extra)\n"); // @[Monitor.scala 255:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_308 & ~_T_1557) begin
          $fatal; // @[Monitor.scala 255:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_316 & ~_T_1329) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries unmanaged address (connected at HellaCache.scala:220:21)\n    at Monitor.scala:259 assert (address_ok, \"'C' channel HintAck carries unmanaged address\" + extra)\n"); // @[Monitor.scala 259:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_316 & ~_T_1329) begin
          $fatal; // @[Monitor.scala 259:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_316 & ~_T_1332) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid source ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:260 assert (source_ok, \"'C' channel HintAck carries invalid source ID\" + extra)\n"); // @[Monitor.scala 260:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_316 & ~_T_1332) begin
          $fatal; // @[Monitor.scala 260:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_316 & ~_T_1339) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck address not aligned to size (connected at HellaCache.scala:220:21)\n    at Monitor.scala:261 assert (is_aligned, \"'C' channel HintAck address not aligned to size\" + extra)\n"); // @[Monitor.scala 261:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_316 & ~_T_1339) begin
          $fatal; // @[Monitor.scala 261:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_316 & ~_T_1557) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid param (connected at HellaCache.scala:220:21)\n    at Monitor.scala:262 assert (bundle.param === UInt(0), \"'C' channel HintAck carries invalid param\" + extra)\n"); // @[Monitor.scala 262:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_316 & ~_T_1557) begin
          $fatal; // @[Monitor.scala 262:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1632 & ~_T_1635) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at HellaCache.scala:220:21)\n    at Monitor.scala:355 assert (a.bits.opcode === opcode, \"'A' channel opcode changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 355:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1632 & ~_T_1635) begin
          $fatal; // @[Monitor.scala 355:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1632 & ~_T_1639) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at HellaCache.scala:220:21)\n    at Monitor.scala:356 assert (a.bits.param  === param,  \"'A' channel param changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 356:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1632 & ~_T_1639) begin
          $fatal; // @[Monitor.scala 356:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1632 & ~_T_1643) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at HellaCache.scala:220:21)\n    at Monitor.scala:357 assert (a.bits.size   === size,   \"'A' channel size changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 357:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1632 & ~_T_1643) begin
          $fatal; // @[Monitor.scala 357:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1632 & ~_T_1647) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at HellaCache.scala:220:21)\n    at Monitor.scala:358 assert (a.bits.source === source, \"'A' channel source changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 358:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1632 & ~_T_1647) begin
          $fatal; // @[Monitor.scala 358:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1632 & ~_T_1651) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at HellaCache.scala:220:21)\n    at Monitor.scala:359 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); // @[Monitor.scala 359:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1632 & ~_T_1651) begin
          $fatal; // @[Monitor.scala 359:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1689 & ~_T_1692) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at HellaCache.scala:220:21)\n    at Monitor.scala:425 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 425:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1689 & ~_T_1692) begin
          $fatal; // @[Monitor.scala 425:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1689 & ~_T_1696) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at HellaCache.scala:220:21)\n    at Monitor.scala:426 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 426:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1689 & ~_T_1696) begin
          $fatal; // @[Monitor.scala 426:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1689 & ~_T_1700) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at HellaCache.scala:220:21)\n    at Monitor.scala:427 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 427:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1689 & ~_T_1700) begin
          $fatal; // @[Monitor.scala 427:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1689 & ~_T_1704) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at HellaCache.scala:220:21)\n    at Monitor.scala:428 assert (d.bits.source === source, \"'D' channel source changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 428:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1689 & ~_T_1704) begin
          $fatal; // @[Monitor.scala 428:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1689 & ~_T_1708) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at HellaCache.scala:220:21)\n    at Monitor.scala:429 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); // @[Monitor.scala 429:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1689 & ~_T_1708) begin
          $fatal; // @[Monitor.scala 429:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1689 & ~_T_1712) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at HellaCache.scala:220:21)\n    at Monitor.scala:430 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); // @[Monitor.scala 430:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1689 & ~_T_1712) begin
          $fatal; // @[Monitor.scala 430:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1749 & ~_T_1752) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel opcode changed within multibeat operation (connected at HellaCache.scala:220:21)\n    at Monitor.scala:378 assert (b.bits.opcode === opcode, \"'B' channel opcode changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 378:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1749 & ~_T_1752) begin
          $fatal; // @[Monitor.scala 378:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1749 & ~_T_1756) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel param changed within multibeat operation (connected at HellaCache.scala:220:21)\n    at Monitor.scala:379 assert (b.bits.param  === param,  \"'B' channel param changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 379:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1749 & ~_T_1756) begin
          $fatal; // @[Monitor.scala 379:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1749 & ~_T_1760) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel size changed within multibeat operation (connected at HellaCache.scala:220:21)\n    at Monitor.scala:380 assert (b.bits.size   === size,   \"'B' channel size changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 380:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1749 & ~_T_1760) begin
          $fatal; // @[Monitor.scala 380:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1749 & ~_T_1764) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel source changed within multibeat operation (connected at HellaCache.scala:220:21)\n    at Monitor.scala:381 assert (b.bits.source === source, \"'B' channel source changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 381:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1749 & ~_T_1764) begin
          $fatal; // @[Monitor.scala 381:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1749 & ~_T_1768) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel addresss changed with multibeat operation (connected at HellaCache.scala:220:21)\n    at Monitor.scala:382 assert (b.bits.address=== address,\"'B' channel addresss changed with multibeat operation\" + extra)\n"); // @[Monitor.scala 382:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1749 & ~_T_1768) begin
          $fatal; // @[Monitor.scala 382:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1804 & ~_T_1807) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel opcode changed within multibeat operation (connected at HellaCache.scala:220:21)\n    at Monitor.scala:401 assert (c.bits.opcode === opcode, \"'C' channel opcode changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 401:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1804 & ~_T_1807) begin
          $fatal; // @[Monitor.scala 401:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1804 & ~_T_1811) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel param changed within multibeat operation (connected at HellaCache.scala:220:21)\n    at Monitor.scala:402 assert (c.bits.param  === param,  \"'C' channel param changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 402:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1804 & ~_T_1811) begin
          $fatal; // @[Monitor.scala 402:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1804 & ~_T_1815) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel size changed within multibeat operation (connected at HellaCache.scala:220:21)\n    at Monitor.scala:403 assert (c.bits.size   === size,   \"'C' channel size changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 403:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1804 & ~_T_1815) begin
          $fatal; // @[Monitor.scala 403:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1804 & ~_T_1819) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel source changed within multibeat operation (connected at HellaCache.scala:220:21)\n    at Monitor.scala:404 assert (c.bits.source === source, \"'C' channel source changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 404:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1804 & ~_T_1819) begin
          $fatal; // @[Monitor.scala 404:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1804 & ~_T_1823) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel address changed with multibeat operation (connected at HellaCache.scala:220:21)\n    at Monitor.scala:405 assert (c.bits.address=== address,\"'C' channel address changed with multibeat operation\" + extra)\n"); // @[Monitor.scala 405:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1804 & ~_T_1823) begin
          $fatal; // @[Monitor.scala 405:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1875 & ~_T_1882) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:460 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); // @[Monitor.scala 460:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1875 & ~_T_1882) begin
          $fatal; // @[Monitor.scala 460:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1891 & ~_T_1897) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at HellaCache.scala:220:21)\n    at Monitor.scala:467 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); // @[Monitor.scala 467:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1891 & ~_T_1897) begin
          $fatal; // @[Monitor.scala 467:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_1904) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at HellaCache.scala:220:21)\n    at Monitor.scala:471 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); // @[Monitor.scala 471:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_1904) begin
          $fatal; // @[Monitor.scala 471:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1956 & ~_T_1962) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel re-used a sink ID (connected at HellaCache.scala:220:21)\n    at Monitor.scala:494 assert(!inflight(bundle.d.bits.sink), \"'D' channel re-used a sink ID\" + extra)\n"); // @[Monitor.scala 494:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1956 & ~_T_1962) begin
          $fatal; // @[Monitor.scala 494:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1966 & ~_T_1974) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel acknowledged for nothing inflight (connected at HellaCache.scala:220:21)\n    at Monitor.scala:500 assert((d_set | inflight)(bundle.e.bits.sink), \"'E' channel acknowledged for nothing inflight\" + extra)\n"); // @[Monitor.scala 500:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1966 & ~_T_1974) begin
          $fatal; // @[Monitor.scala 500:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    if (metaReset) begin
      TLMonitor_64_metaAssert <= 1'h0;
    end else begin
      TLMonitor_64_metaAssert <= TLMonitor_64_metaAssert | TLMonitor_64_or0;
    end
  end
endmodule
module TLMonitor_65(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [31:0] io_in_a_bits_address,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [1:0]  io_in_d_bits_param,
  input  [3:0]  io_in_d_bits_size,
  input  [1:0]  io_in_d_bits_sink,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [31:0] _T_32; // @[Edges.scala 21:16]
  wire  _T_33; // @[Edges.scala 21:24]
  wire [32:0] _T_101; // @[Parameters.scala 121:49]
  wire [31:0] _T_114; // @[Parameters.scala 121:31]
  wire [32:0] _T_115; // @[Parameters.scala 121:49]
  wire [32:0] _T_117; // @[Parameters.scala 121:52]
  wire  _T_118; // @[Parameters.scala 121:67]
  wire [31:0] _T_121; // @[Parameters.scala 121:31]
  wire [32:0] _T_122; // @[Parameters.scala 121:49]
  wire [32:0] _T_124; // @[Parameters.scala 121:52]
  wire  _T_125; // @[Parameters.scala 121:67]
  wire [31:0] _T_126; // @[Parameters.scala 121:31]
  wire [32:0] _T_127; // @[Parameters.scala 121:49]
  wire [32:0] _T_129; // @[Parameters.scala 121:52]
  wire  _T_130; // @[Parameters.scala 121:67]
  wire [31:0] _T_131; // @[Parameters.scala 121:31]
  wire [32:0] _T_132; // @[Parameters.scala 121:49]
  wire [32:0] _T_134; // @[Parameters.scala 121:52]
  wire  _T_135; // @[Parameters.scala 121:67]
  wire [32:0] _T_139; // @[Parameters.scala 121:52]
  wire  _T_140; // @[Parameters.scala 121:67]
  wire [31:0] _T_141; // @[Parameters.scala 121:31]
  wire [32:0] _T_142; // @[Parameters.scala 121:49]
  wire [32:0] _T_144; // @[Parameters.scala 121:52]
  wire  _T_145; // @[Parameters.scala 121:67]
  wire [31:0] _T_146; // @[Parameters.scala 121:31]
  wire [32:0] _T_147; // @[Parameters.scala 121:49]
  wire [32:0] _T_149; // @[Parameters.scala 121:52]
  wire  _T_150; // @[Parameters.scala 121:67]
  wire  _T_173; // @[Monitor.scala 53:14]
  wire  _T_316; // @[Parameters.scala 169:42]
  wire  _T_317; // @[Parameters.scala 169:42]
  wire  _T_318; // @[Parameters.scala 169:42]
  wire  _T_319; // @[Parameters.scala 169:42]
  wire  _T_320; // @[Parameters.scala 169:42]
  wire  _T_323; // @[Parameters.scala 170:30]
  wire  _T_325; // @[Monitor.scala 72:14]
  wire  _T_702; // @[Bundles.scala 43:24]
  wire  _T_704; // @[Monitor.scala 268:12]
  wire  _T_715; // @[Monitor.scala 275:25]
  wire  _T_719; // @[Monitor.scala 277:27]
  wire  _T_721; // @[Monitor.scala 277:14]
  wire  _T_723; // @[Monitor.scala 278:28]
  wire  _T_725; // @[Monitor.scala 278:14]
  wire  _T_729; // @[Monitor.scala 279:14]
  wire  _T_733; // @[Monitor.scala 280:14]
  wire  _T_735; // @[Monitor.scala 283:25]
  wire  _T_746; // @[Bundles.scala 103:26]
  wire  _T_748; // @[Monitor.scala 287:14]
  wire  _T_750; // @[Monitor.scala 288:28]
  wire  _T_752; // @[Monitor.scala 288:14]
  wire  _T_763; // @[Monitor.scala 293:25]
  wire  _T_783; // @[Monitor.scala 299:30]
  wire  _T_785; // @[Monitor.scala 299:14]
  wire  _T_792; // @[Monitor.scala 303:25]
  wire  _T_809; // @[Monitor.scala 311:25]
  wire  _T_827; // @[Monitor.scala 319:25]
  wire  _T_856; // @[Bundles.scala 277:22]
  reg [8:0] _T_866; // @[Edges.scala 229:27]
  reg [31:0] _RAND_0;
  wire [8:0] _T_869; // @[Edges.scala 230:28]
  wire  _T_870; // @[Edges.scala 231:25]
  reg [31:0] _T_887; // @[Monitor.scala 353:22]
  reg [31:0] _RAND_1;
  wire  _T_889; // @[Monitor.scala 354:19]
  wire  _T_906; // @[Monitor.scala 359:29]
  wire  _T_908; // @[Monitor.scala 359:14]
  wire  _T_911; // @[Monitor.scala 361:20]
  wire [26:0] _T_914; // @[package.scala 185:77]
  wire [8:0] _T_917; // @[Edges.scala 220:59]
  reg [8:0] _T_921; // @[Edges.scala 229:27]
  reg [31:0] _RAND_2;
  wire [8:0] _T_924; // @[Edges.scala 230:28]
  wire  _T_925; // @[Edges.scala 231:25]
  reg [2:0] _T_934; // @[Monitor.scala 418:22]
  reg [31:0] _RAND_3;
  reg [1:0] _T_936; // @[Monitor.scala 419:22]
  reg [31:0] _RAND_4;
  reg [3:0] _T_938; // @[Monitor.scala 420:22]
  reg [31:0] _RAND_5;
  reg [1:0] _T_942; // @[Monitor.scala 422:22]
  reg [31:0] _RAND_6;
  reg  _T_944; // @[Monitor.scala 423:22]
  reg [31:0] _RAND_7;
  wire  _T_946; // @[Monitor.scala 424:19]
  wire  _T_947; // @[Monitor.scala 425:29]
  wire  _T_949; // @[Monitor.scala 425:14]
  wire  _T_951; // @[Monitor.scala 426:29]
  wire  _T_953; // @[Monitor.scala 426:14]
  wire  _T_955; // @[Monitor.scala 427:29]
  wire  _T_957; // @[Monitor.scala 427:14]
  wire  _T_963; // @[Monitor.scala 429:29]
  wire  _T_965; // @[Monitor.scala 429:14]
  wire  _T_967; // @[Monitor.scala 430:29]
  wire  _T_969; // @[Monitor.scala 430:14]
  wire  _T_972; // @[Monitor.scala 432:20]
  reg  _T_974; // @[Monitor.scala 452:27]
  reg [31:0] _RAND_8;
  reg [8:0] _T_985; // @[Edges.scala 229:27]
  reg [31:0] _RAND_9;
  wire [8:0] _T_988; // @[Edges.scala 230:28]
  wire  _T_989; // @[Edges.scala 231:25]
  reg [8:0] _T_1006; // @[Edges.scala 229:27]
  reg [31:0] _RAND_10;
  wire [8:0] _T_1009; // @[Edges.scala 230:28]
  wire  _T_1010; // @[Edges.scala 231:25]
  wire  _T_1021; // @[Monitor.scala 458:27]
  wire  _T_1028; // @[Monitor.scala 460:13]
  wire [1:0] _GEN_15; // @[Monitor.scala 458:72]
  wire  _T_1034; // @[Monitor.scala 465:27]
  wire  _T_1037; // @[Monitor.scala 465:72]
  wire  _T_1039; // @[Monitor.scala 467:21]
  wire  _T_1043; // @[Monitor.scala 467:13]
  wire [1:0] _GEN_16; // @[Monitor.scala 465:91]
  wire  _T_1045; // @[Monitor.scala 471:20]
  wire  _T_1048; // @[Monitor.scala 471:30]
  wire  _T_1050; // @[Monitor.scala 471:13]
  wire  _T_1052; // @[Monitor.scala 474:27]
  wire  _T_1054; // @[Monitor.scala 474:36]
  wire  _GEN_18; // @[Monitor.scala 277:14]
  wire  _GEN_26; // @[Monitor.scala 286:14]
  wire  _GEN_34; // @[Monitor.scala 296:14]
  wire  _GEN_42; // @[Monitor.scala 306:14]
  wire  _GEN_46; // @[Monitor.scala 314:14]
  wire  _GEN_50; // @[Monitor.scala 322:14]
  wire [29:0] TLMonitor_65_covSum;
  wire  stopEn0;
  wire  stopEn1;
  wire  stopEn2;
  wire  stopEn3;
  wire  stopEn4;
  wire  stopEn5;
  wire  stopEn6;
  wire  stopEn7;
  wire  stopEn8;
  wire  stopEn9;
  wire  stopEn10;
  wire  stopEn11;
  wire  stopEn12;
  wire  stopEn13;
  wire  stopEn14;
  wire  stopEn15;
  wire  stopEn16;
  wire  stopEn17;
  wire  stopEn18;
  wire  stopEn19;
  wire  stopEn20;
  wire  stopEn21;
  wire  stopEn22;
  wire  stopEn23;
  wire  stopEn24;
  wire  stopEn25;
  wire  stopEn26;
  wire  stopEn27;
  wire  stopEn28;
  wire  stopEn29;
  wire  TLMonitor_65_or16;
  wire  TLMonitor_65_or7;
  wire  TLMonitor_65_or17;
  wire  TLMonitor_65_or18;
  wire  TLMonitor_65_or8;
  wire  TLMonitor_65_or3;
  wire  TLMonitor_65_or19;
  wire  TLMonitor_65_or20;
  wire  TLMonitor_65_or9;
  wire  TLMonitor_65_or21;
  wire  TLMonitor_65_or22;
  wire  TLMonitor_65_or10;
  wire  TLMonitor_65_or4;
  wire  TLMonitor_65_or1;
  wire  TLMonitor_65_or24;
  wire  TLMonitor_65_or11;
  wire  TLMonitor_65_or25;
  wire  TLMonitor_65_or26;
  wire  TLMonitor_65_or12;
  wire  TLMonitor_65_or5;
  wire  TLMonitor_65_or27;
  wire  TLMonitor_65_or28;
  wire  TLMonitor_65_or13;
  wire  TLMonitor_65_or29;
  wire  TLMonitor_65_or30;
  wire  TLMonitor_65_or14;
  wire  TLMonitor_65_or6;
  wire  TLMonitor_65_or2;
  wire  TLMonitor_65_or0;
  reg  TLMonitor_65_metaAssert;
  reg [31:0] _RAND_11;
  assign _T_32 = io_in_a_bits_address & 32'h3f; // @[Edges.scala 21:16]
  assign _T_33 = _T_32 == 32'h0; // @[Edges.scala 21:24]
  assign _T_101 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 121:49]
  assign _T_114 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 121:31]
  assign _T_115 = {1'b0,$signed(_T_114)}; // @[Parameters.scala 121:49]
  assign _T_117 = $signed(_T_115) & -33'sh10000000; // @[Parameters.scala 121:52]
  assign _T_118 = $signed(_T_117) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_121 = io_in_a_bits_address ^ 32'h3000; // @[Parameters.scala 121:31]
  assign _T_122 = {1'b0,$signed(_T_121)}; // @[Parameters.scala 121:49]
  assign _T_124 = $signed(_T_122) & -33'sh1000; // @[Parameters.scala 121:52]
  assign _T_125 = $signed(_T_124) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_126 = io_in_a_bits_address ^ 32'hc000000; // @[Parameters.scala 121:31]
  assign _T_127 = {1'b0,$signed(_T_126)}; // @[Parameters.scala 121:49]
  assign _T_129 = $signed(_T_127) & -33'sh4000000; // @[Parameters.scala 121:52]
  assign _T_130 = $signed(_T_129) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_131 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 121:31]
  assign _T_132 = {1'b0,$signed(_T_131)}; // @[Parameters.scala 121:49]
  assign _T_134 = $signed(_T_132) & -33'sh10000; // @[Parameters.scala 121:52]
  assign _T_135 = $signed(_T_134) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_139 = $signed(_T_101) & -33'sh1000; // @[Parameters.scala 121:52]
  assign _T_140 = $signed(_T_139) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_141 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 121:31]
  assign _T_142 = {1'b0,$signed(_T_141)}; // @[Parameters.scala 121:49]
  assign _T_144 = $signed(_T_142) & -33'sh10000; // @[Parameters.scala 121:52]
  assign _T_145 = $signed(_T_144) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_146 = io_in_a_bits_address ^ 32'h60000000; // @[Parameters.scala 121:31]
  assign _T_147 = {1'b0,$signed(_T_146)}; // @[Parameters.scala 121:49]
  assign _T_149 = $signed(_T_147) & -33'sh20000000; // @[Parameters.scala 121:52]
  assign _T_150 = $signed(_T_149) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_173 = _T_33 | reset; // @[Monitor.scala 53:14]
  assign _T_316 = _T_130 | _T_135; // @[Parameters.scala 169:42]
  assign _T_317 = _T_316 | _T_140; // @[Parameters.scala 169:42]
  assign _T_318 = _T_317 | _T_145; // @[Parameters.scala 169:42]
  assign _T_319 = _T_318 | _T_118; // @[Parameters.scala 169:42]
  assign _T_320 = _T_319 | _T_150; // @[Parameters.scala 169:42]
  assign _T_323 = _T_125 | _T_320; // @[Parameters.scala 170:30]
  assign _T_325 = _T_323 | reset; // @[Monitor.scala 72:14]
  assign _T_702 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 43:24]
  assign _T_704 = _T_702 | reset; // @[Monitor.scala 268:12]
  assign _T_715 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 275:25]
  assign _T_719 = io_in_d_bits_size >= 4'h3; // @[Monitor.scala 277:27]
  assign _T_721 = _T_719 | reset; // @[Monitor.scala 277:14]
  assign _T_723 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 278:28]
  assign _T_725 = _T_723 | reset; // @[Monitor.scala 278:14]
  assign _T_729 = ~io_in_d_bits_corrupt | reset; // @[Monitor.scala 279:14]
  assign _T_733 = ~io_in_d_bits_denied | reset; // @[Monitor.scala 280:14]
  assign _T_735 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 283:25]
  assign _T_746 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 103:26]
  assign _T_748 = _T_746 | reset; // @[Monitor.scala 287:14]
  assign _T_750 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 288:28]
  assign _T_752 = _T_750 | reset; // @[Monitor.scala 288:14]
  assign _T_763 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 293:25]
  assign _T_783 = ~io_in_d_bits_denied | io_in_d_bits_corrupt; // @[Monitor.scala 299:30]
  assign _T_785 = _T_783 | reset; // @[Monitor.scala 299:14]
  assign _T_792 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 303:25]
  assign _T_809 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 311:25]
  assign _T_827 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 319:25]
  assign _T_856 = io_in_a_ready & io_in_a_valid; // @[Bundles.scala 277:22]
  assign _T_869 = _T_866 - 9'h1; // @[Edges.scala 230:28]
  assign _T_870 = _T_866 == 9'h0; // @[Edges.scala 231:25]
  assign _T_889 = io_in_a_valid & ~_T_870; // @[Monitor.scala 354:19]
  assign _T_906 = io_in_a_bits_address == _T_887; // @[Monitor.scala 359:29]
  assign _T_908 = _T_906 | reset; // @[Monitor.scala 359:14]
  assign _T_911 = _T_856 & _T_870; // @[Monitor.scala 361:20]
  assign _T_914 = 27'hfff << io_in_d_bits_size; // @[package.scala 185:77]
  assign _T_917 = ~_T_914[11:3]; // @[Edges.scala 220:59]
  assign _T_924 = _T_921 - 9'h1; // @[Edges.scala 230:28]
  assign _T_925 = _T_921 == 9'h0; // @[Edges.scala 231:25]
  assign _T_946 = io_in_d_valid & ~_T_925; // @[Monitor.scala 424:19]
  assign _T_947 = io_in_d_bits_opcode == _T_934; // @[Monitor.scala 425:29]
  assign _T_949 = _T_947 | reset; // @[Monitor.scala 425:14]
  assign _T_951 = io_in_d_bits_param == _T_936; // @[Monitor.scala 426:29]
  assign _T_953 = _T_951 | reset; // @[Monitor.scala 426:14]
  assign _T_955 = io_in_d_bits_size == _T_938; // @[Monitor.scala 427:29]
  assign _T_957 = _T_955 | reset; // @[Monitor.scala 427:14]
  assign _T_963 = io_in_d_bits_sink == _T_942; // @[Monitor.scala 429:29]
  assign _T_965 = _T_963 | reset; // @[Monitor.scala 429:14]
  assign _T_967 = io_in_d_bits_denied == _T_944; // @[Monitor.scala 430:29]
  assign _T_969 = _T_967 | reset; // @[Monitor.scala 430:14]
  assign _T_972 = io_in_d_valid & _T_925; // @[Monitor.scala 432:20]
  assign _T_988 = _T_985 - 9'h1; // @[Edges.scala 230:28]
  assign _T_989 = _T_985 == 9'h0; // @[Edges.scala 231:25]
  assign _T_1009 = _T_1006 - 9'h1; // @[Edges.scala 230:28]
  assign _T_1010 = _T_1006 == 9'h0; // @[Edges.scala 231:25]
  assign _T_1021 = _T_856 & _T_989; // @[Monitor.scala 458:27]
  assign _T_1028 = ~_T_974 | reset; // @[Monitor.scala 460:13]
  assign _GEN_15 = _T_1021 ? 2'h1 : 2'h0; // @[Monitor.scala 458:72]
  assign _T_1034 = io_in_d_valid & _T_1010; // @[Monitor.scala 465:27]
  assign _T_1037 = _T_1034 & ~_T_715; // @[Monitor.scala 465:72]
  assign _T_1039 = _GEN_15[0] | _T_974; // @[Monitor.scala 467:21]
  assign _T_1043 = _T_1039 | reset; // @[Monitor.scala 467:13]
  assign _GEN_16 = _T_1037 ? 2'h1 : 2'h0; // @[Monitor.scala 465:91]
  assign _T_1045 = _GEN_15[0] != _GEN_16[0]; // @[Monitor.scala 471:20]
  assign _T_1048 = _T_1045 | ~_GEN_15[0]; // @[Monitor.scala 471:30]
  assign _T_1050 = _T_1048 | reset; // @[Monitor.scala 471:13]
  assign _T_1052 = _T_974 | _GEN_15[0]; // @[Monitor.scala 474:27]
  assign _T_1054 = _T_1052 & ~_GEN_16[0]; // @[Monitor.scala 474:36]
  assign _GEN_18 = io_in_d_valid & _T_715; // @[Monitor.scala 277:14]
  assign _GEN_26 = io_in_d_valid & _T_735; // @[Monitor.scala 286:14]
  assign _GEN_34 = io_in_d_valid & _T_763; // @[Monitor.scala 296:14]
  assign _GEN_42 = io_in_d_valid & _T_792; // @[Monitor.scala 306:14]
  assign _GEN_46 = io_in_d_valid & _T_809; // @[Monitor.scala 314:14]
  assign _GEN_50 = io_in_d_valid & _T_827; // @[Monitor.scala 322:14]
  assign TLMonitor_65_covSum = 30'h0;
  assign io_covSum = TLMonitor_65_covSum;
  assign stopEn0 = io_in_a_valid & ~_T_325;
  assign stopEn1 = io_in_a_valid & ~_T_173;
  assign stopEn2 = io_in_d_valid & ~_T_704;
  assign stopEn3 = _GEN_18 & ~_T_721;
  assign stopEn4 = _GEN_18 & ~_T_725;
  assign stopEn5 = _GEN_18 & ~_T_729;
  assign stopEn6 = _GEN_18 & ~_T_733;
  assign stopEn7 = _GEN_26 & ~_T_721;
  assign stopEn8 = _GEN_26 & ~_T_748;
  assign stopEn9 = _GEN_26 & ~_T_752;
  assign stopEn10 = _GEN_26 & ~_T_729;
  assign stopEn11 = _GEN_34 & ~_T_721;
  assign stopEn12 = _GEN_34 & ~_T_748;
  assign stopEn13 = _GEN_34 & ~_T_752;
  assign stopEn14 = _GEN_34 & ~_T_785;
  assign stopEn15 = _GEN_42 & ~_T_725;
  assign stopEn16 = _GEN_42 & ~_T_729;
  assign stopEn17 = _GEN_46 & ~_T_725;
  assign stopEn18 = _GEN_46 & ~_T_785;
  assign stopEn19 = _GEN_50 & ~_T_725;
  assign stopEn20 = _GEN_50 & ~_T_729;
  assign stopEn21 = _T_889 & ~_T_908;
  assign stopEn22 = _T_946 & ~_T_949;
  assign stopEn23 = _T_946 & ~_T_953;
  assign stopEn24 = _T_946 & ~_T_957;
  assign stopEn25 = _T_946 & ~_T_965;
  assign stopEn26 = _T_946 & ~_T_969;
  assign stopEn27 = _T_1021 & ~_T_1028;
  assign stopEn28 = _T_1037 & ~_T_1043;
  assign stopEn29 = ~_T_1050;
  assign TLMonitor_65_or16 = stopEn1 | stopEn2;
  assign TLMonitor_65_or7 = stopEn0 | TLMonitor_65_or16;
  assign TLMonitor_65_or17 = stopEn3 | stopEn4;
  assign TLMonitor_65_or18 = stopEn5 | stopEn6;
  assign TLMonitor_65_or8 = TLMonitor_65_or17 | TLMonitor_65_or18;
  assign TLMonitor_65_or3 = TLMonitor_65_or7 | TLMonitor_65_or8;
  assign TLMonitor_65_or19 = stopEn7 | stopEn8;
  assign TLMonitor_65_or20 = stopEn9 | stopEn10;
  assign TLMonitor_65_or9 = TLMonitor_65_or19 | TLMonitor_65_or20;
  assign TLMonitor_65_or21 = stopEn11 | stopEn12;
  assign TLMonitor_65_or22 = stopEn13 | stopEn14;
  assign TLMonitor_65_or10 = TLMonitor_65_or21 | TLMonitor_65_or22;
  assign TLMonitor_65_or4 = TLMonitor_65_or9 | TLMonitor_65_or10;
  assign TLMonitor_65_or1 = TLMonitor_65_or3 | TLMonitor_65_or4;
  assign TLMonitor_65_or24 = stopEn16 | stopEn17;
  assign TLMonitor_65_or11 = stopEn15 | TLMonitor_65_or24;
  assign TLMonitor_65_or25 = stopEn18 | stopEn19;
  assign TLMonitor_65_or26 = stopEn20 | stopEn21;
  assign TLMonitor_65_or12 = TLMonitor_65_or25 | TLMonitor_65_or26;
  assign TLMonitor_65_or5 = TLMonitor_65_or11 | TLMonitor_65_or12;
  assign TLMonitor_65_or27 = stopEn22 | stopEn23;
  assign TLMonitor_65_or28 = stopEn24 | stopEn25;
  assign TLMonitor_65_or13 = TLMonitor_65_or27 | TLMonitor_65_or28;
  assign TLMonitor_65_or29 = stopEn26 | stopEn27;
  assign TLMonitor_65_or30 = stopEn28 | stopEn29;
  assign TLMonitor_65_or14 = TLMonitor_65_or29 | TLMonitor_65_or30;
  assign TLMonitor_65_or6 = TLMonitor_65_or13 | TLMonitor_65_or14;
  assign TLMonitor_65_or2 = TLMonitor_65_or5 | TLMonitor_65_or6;
  assign TLMonitor_65_or0 = TLMonitor_65_or1 | TLMonitor_65_or2;
  assign metaAssert = TLMonitor_65_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_866 = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_887 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_921 = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_934 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_936 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_938 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_942 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_944 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_974 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_985 = _RAND_9[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_1006 = _RAND_10[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  TLMonitor_65_metaAssert = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      _T_866 <= 9'h0;
    end else if (reset) begin
      _T_866 <= 9'h0;
    end else if (_T_856) begin
      if (_T_870) begin
        _T_866 <= 9'h0;
      end else begin
        _T_866 <= _T_869;
      end
    end
    if (metaReset) begin
      _T_887 <= 32'h0;
    end else if (_T_911) begin
      _T_887 <= io_in_a_bits_address;
    end
    if (metaReset) begin
      _T_921 <= 9'h0;
    end else if (reset) begin
      _T_921 <= 9'h0;
    end else if (io_in_d_valid) begin
      if (_T_925) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_921 <= _T_917;
        end else begin
          _T_921 <= 9'h0;
        end
      end else begin
        _T_921 <= _T_924;
      end
    end
    if (metaReset) begin
      _T_934 <= 3'h0;
    end else if (_T_972) begin
      _T_934 <= io_in_d_bits_opcode;
    end
    if (metaReset) begin
      _T_936 <= 2'h0;
    end else if (_T_972) begin
      _T_936 <= io_in_d_bits_param;
    end
    if (metaReset) begin
      _T_938 <= 4'h0;
    end else if (_T_972) begin
      _T_938 <= io_in_d_bits_size;
    end
    if (metaReset) begin
      _T_942 <= 2'h0;
    end else if (_T_972) begin
      _T_942 <= io_in_d_bits_sink;
    end
    if (metaReset) begin
      _T_944 <= 1'h0;
    end else if (_T_972) begin
      _T_944 <= io_in_d_bits_denied;
    end
    if (metaReset) begin
      _T_974 <= 1'h0;
    end else if (reset) begin
      _T_974 <= 1'h0;
    end else begin
      _T_974 <= _T_1054;
    end
    if (metaReset) begin
      _T_985 <= 9'h0;
    end else if (reset) begin
      _T_985 <= 9'h0;
    end else if (_T_856) begin
      if (_T_989) begin
        _T_985 <= 9'h0;
      end else begin
        _T_985 <= _T_988;
      end
    end
    if (metaReset) begin
      _T_1006 <= 9'h0;
    end else if (reset) begin
      _T_1006 <= 9'h0;
    end else if (io_in_d_valid) begin
      if (_T_1010) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1006 <= _T_917;
        end else begin
          _T_1006 <= 9'h0;
        end
      end else begin
        _T_1006 <= _T_1009;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & ~_T_325) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at Frontend.scala:341:21)\n    at Monitor.scala:72 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); // @[Monitor.scala 72:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & ~_T_325) begin
          $fatal; // @[Monitor.scala 72:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & ~_T_173) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at Frontend.scala:341:21)\n    at Monitor.scala:74 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); // @[Monitor.scala 74:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & ~_T_173) begin
          $fatal; // @[Monitor.scala 74:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~_T_704) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at Frontend.scala:341:21)\n    at Monitor.scala:268 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); // @[Monitor.scala 268:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~_T_704) begin
          $fatal; // @[Monitor.scala 268:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_18 & ~_T_721) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at Frontend.scala:341:21)\n    at Monitor.scala:277 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); // @[Monitor.scala 277:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_18 & ~_T_721) begin
          $fatal; // @[Monitor.scala 277:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_18 & ~_T_725) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at Frontend.scala:341:21)\n    at Monitor.scala:278 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); // @[Monitor.scala 278:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_18 & ~_T_725) begin
          $fatal; // @[Monitor.scala 278:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_18 & ~_T_729) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at Frontend.scala:341:21)\n    at Monitor.scala:279 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); // @[Monitor.scala 279:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_18 & ~_T_729) begin
          $fatal; // @[Monitor.scala 279:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_18 & ~_T_733) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at Frontend.scala:341:21)\n    at Monitor.scala:280 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); // @[Monitor.scala 280:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_18 & ~_T_733) begin
          $fatal; // @[Monitor.scala 280:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_26 & ~_T_721) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at Frontend.scala:341:21)\n    at Monitor.scala:286 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); // @[Monitor.scala 286:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_26 & ~_T_721) begin
          $fatal; // @[Monitor.scala 286:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_26 & ~_T_748) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at Frontend.scala:341:21)\n    at Monitor.scala:287 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); // @[Monitor.scala 287:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_26 & ~_T_748) begin
          $fatal; // @[Monitor.scala 287:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_26 & ~_T_752) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at Frontend.scala:341:21)\n    at Monitor.scala:288 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); // @[Monitor.scala 288:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_26 & ~_T_752) begin
          $fatal; // @[Monitor.scala 288:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_26 & ~_T_729) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at Frontend.scala:341:21)\n    at Monitor.scala:289 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); // @[Monitor.scala 289:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_26 & ~_T_729) begin
          $fatal; // @[Monitor.scala 289:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_34 & ~_T_721) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at Frontend.scala:341:21)\n    at Monitor.scala:296 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); // @[Monitor.scala 296:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_34 & ~_T_721) begin
          $fatal; // @[Monitor.scala 296:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_34 & ~_T_748) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at Frontend.scala:341:21)\n    at Monitor.scala:297 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); // @[Monitor.scala 297:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_34 & ~_T_748) begin
          $fatal; // @[Monitor.scala 297:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_34 & ~_T_752) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at Frontend.scala:341:21)\n    at Monitor.scala:298 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); // @[Monitor.scala 298:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_34 & ~_T_752) begin
          $fatal; // @[Monitor.scala 298:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_34 & ~_T_785) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at Frontend.scala:341:21)\n    at Monitor.scala:299 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); // @[Monitor.scala 299:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_34 & ~_T_785) begin
          $fatal; // @[Monitor.scala 299:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_42 & ~_T_725) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at Frontend.scala:341:21)\n    at Monitor.scala:306 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); // @[Monitor.scala 306:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_42 & ~_T_725) begin
          $fatal; // @[Monitor.scala 306:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_42 & ~_T_729) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at Frontend.scala:341:21)\n    at Monitor.scala:307 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); // @[Monitor.scala 307:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_42 & ~_T_729) begin
          $fatal; // @[Monitor.scala 307:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_46 & ~_T_725) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at Frontend.scala:341:21)\n    at Monitor.scala:314 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); // @[Monitor.scala 314:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_46 & ~_T_725) begin
          $fatal; // @[Monitor.scala 314:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_46 & ~_T_785) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at Frontend.scala:341:21)\n    at Monitor.scala:315 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); // @[Monitor.scala 315:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_46 & ~_T_785) begin
          $fatal; // @[Monitor.scala 315:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_50 & ~_T_725) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at Frontend.scala:341:21)\n    at Monitor.scala:322 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); // @[Monitor.scala 322:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_50 & ~_T_725) begin
          $fatal; // @[Monitor.scala 322:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_50 & ~_T_729) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at Frontend.scala:341:21)\n    at Monitor.scala:323 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); // @[Monitor.scala 323:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_50 & ~_T_729) begin
          $fatal; // @[Monitor.scala 323:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_889 & ~_T_908) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at Frontend.scala:341:21)\n    at Monitor.scala:359 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); // @[Monitor.scala 359:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_889 & ~_T_908) begin
          $fatal; // @[Monitor.scala 359:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_946 & ~_T_949) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at Frontend.scala:341:21)\n    at Monitor.scala:425 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 425:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_946 & ~_T_949) begin
          $fatal; // @[Monitor.scala 425:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_946 & ~_T_953) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at Frontend.scala:341:21)\n    at Monitor.scala:426 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 426:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_946 & ~_T_953) begin
          $fatal; // @[Monitor.scala 426:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_946 & ~_T_957) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at Frontend.scala:341:21)\n    at Monitor.scala:427 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 427:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_946 & ~_T_957) begin
          $fatal; // @[Monitor.scala 427:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_946 & ~_T_965) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at Frontend.scala:341:21)\n    at Monitor.scala:429 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); // @[Monitor.scala 429:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_946 & ~_T_965) begin
          $fatal; // @[Monitor.scala 429:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_946 & ~_T_969) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at Frontend.scala:341:21)\n    at Monitor.scala:430 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); // @[Monitor.scala 430:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_946 & ~_T_969) begin
          $fatal; // @[Monitor.scala 430:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1021 & ~_T_1028) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at Frontend.scala:341:21)\n    at Monitor.scala:460 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); // @[Monitor.scala 460:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1021 & ~_T_1028) begin
          $fatal; // @[Monitor.scala 460:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1037 & ~_T_1043) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at Frontend.scala:341:21)\n    at Monitor.scala:467 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); // @[Monitor.scala 467:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1037 & ~_T_1043) begin
          $fatal; // @[Monitor.scala 467:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_1050) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at Frontend.scala:341:21)\n    at Monitor.scala:471 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); // @[Monitor.scala 471:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_1050) begin
          $fatal; // @[Monitor.scala 471:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    if (metaReset) begin
      TLMonitor_65_metaAssert <= 1'h0;
    end else begin
      TLMonitor_65_metaAssert <= TLMonitor_65_metaAssert | TLMonitor_65_or0;
    end
  end
endmodule
module Arbiter(
  input         io_in_0_valid,
  input  [39:0] io_in_0_bits_addr,
  input  [5:0]  io_in_0_bits_idx,
  input  [21:0] io_in_0_bits_data,
  input         io_in_2_valid,
  input  [39:0] io_in_2_bits_addr,
  input  [5:0]  io_in_2_bits_idx,
  input  [3:0]  io_in_2_bits_way_en,
  input  [21:0] io_in_2_bits_data,
  input         io_in_3_valid,
  input  [39:0] io_in_3_bits_addr,
  input  [5:0]  io_in_3_bits_idx,
  input  [3:0]  io_in_3_bits_way_en,
  input  [21:0] io_in_3_bits_data,
  output        io_in_4_ready,
  input         io_in_4_valid,
  input  [39:0] io_in_4_bits_addr,
  input  [5:0]  io_in_4_bits_idx,
  input  [3:0]  io_in_4_bits_way_en,
  input  [21:0] io_in_4_bits_data,
  output        io_in_5_ready,
  input         io_in_5_valid,
  input  [39:0] io_in_5_bits_addr,
  input  [5:0]  io_in_5_bits_idx,
  input  [3:0]  io_in_5_bits_way_en,
  input  [21:0] io_in_5_bits_data,
  output        io_in_6_ready,
  input         io_in_6_valid,
  input  [39:0] io_in_6_bits_addr,
  input  [5:0]  io_in_6_bits_idx,
  input  [3:0]  io_in_6_bits_way_en,
  input  [21:0] io_in_6_bits_data,
  output        io_in_7_ready,
  input         io_in_7_valid,
  input  [39:0] io_in_7_bits_addr,
  input  [5:0]  io_in_7_bits_idx,
  input  [3:0]  io_in_7_bits_way_en,
  input  [21:0] io_in_7_bits_data,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_write,
  output [39:0] io_out_bits_addr,
  output [5:0]  io_out_bits_idx,
  output [3:0]  io_out_bits_way_en,
  output [21:0] io_out_bits_data,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [21:0] _GEN_1; // @[Arbiter.scala 126:27]
  wire [3:0] _GEN_2; // @[Arbiter.scala 126:27]
  wire [5:0] _GEN_3; // @[Arbiter.scala 126:27]
  wire [39:0] _GEN_4; // @[Arbiter.scala 126:27]
  wire [21:0] _GEN_7; // @[Arbiter.scala 126:27]
  wire [3:0] _GEN_8; // @[Arbiter.scala 126:27]
  wire [5:0] _GEN_9; // @[Arbiter.scala 126:27]
  wire [39:0] _GEN_10; // @[Arbiter.scala 126:27]
  wire [21:0] _GEN_13; // @[Arbiter.scala 126:27]
  wire [3:0] _GEN_14; // @[Arbiter.scala 126:27]
  wire [5:0] _GEN_15; // @[Arbiter.scala 126:27]
  wire [39:0] _GEN_16; // @[Arbiter.scala 126:27]
  wire [21:0] _GEN_19; // @[Arbiter.scala 126:27]
  wire [3:0] _GEN_20; // @[Arbiter.scala 126:27]
  wire [5:0] _GEN_21; // @[Arbiter.scala 126:27]
  wire [39:0] _GEN_22; // @[Arbiter.scala 126:27]
  wire  _GEN_23; // @[Arbiter.scala 126:27]
  wire [21:0] _GEN_25; // @[Arbiter.scala 126:27]
  wire [3:0] _GEN_26; // @[Arbiter.scala 126:27]
  wire [5:0] _GEN_27; // @[Arbiter.scala 126:27]
  wire [39:0] _GEN_28; // @[Arbiter.scala 126:27]
  wire  _GEN_29; // @[Arbiter.scala 126:27]
  wire  _T_210; // @[Arbiter.scala 31:68]
  wire  _T_211; // @[Arbiter.scala 31:68]
  wire  _T_212; // @[Arbiter.scala 31:68]
  wire  _T_213; // @[Arbiter.scala 31:68]
  wire  _T_214; // @[Arbiter.scala 31:68]
  wire [29:0] Arbiter_covSum;
  assign _GEN_1 = io_in_6_valid ? io_in_6_bits_data : io_in_7_bits_data; // @[Arbiter.scala 126:27]
  assign _GEN_2 = io_in_6_valid ? io_in_6_bits_way_en : io_in_7_bits_way_en; // @[Arbiter.scala 126:27]
  assign _GEN_3 = io_in_6_valid ? io_in_6_bits_idx : io_in_7_bits_idx; // @[Arbiter.scala 126:27]
  assign _GEN_4 = io_in_6_valid ? io_in_6_bits_addr : io_in_7_bits_addr; // @[Arbiter.scala 126:27]
  assign _GEN_7 = io_in_5_valid ? io_in_5_bits_data : _GEN_1; // @[Arbiter.scala 126:27]
  assign _GEN_8 = io_in_5_valid ? io_in_5_bits_way_en : _GEN_2; // @[Arbiter.scala 126:27]
  assign _GEN_9 = io_in_5_valid ? io_in_5_bits_idx : _GEN_3; // @[Arbiter.scala 126:27]
  assign _GEN_10 = io_in_5_valid ? io_in_5_bits_addr : _GEN_4; // @[Arbiter.scala 126:27]
  assign _GEN_13 = io_in_4_valid ? io_in_4_bits_data : _GEN_7; // @[Arbiter.scala 126:27]
  assign _GEN_14 = io_in_4_valid ? io_in_4_bits_way_en : _GEN_8; // @[Arbiter.scala 126:27]
  assign _GEN_15 = io_in_4_valid ? io_in_4_bits_idx : _GEN_9; // @[Arbiter.scala 126:27]
  assign _GEN_16 = io_in_4_valid ? io_in_4_bits_addr : _GEN_10; // @[Arbiter.scala 126:27]
  assign _GEN_19 = io_in_3_valid ? io_in_3_bits_data : _GEN_13; // @[Arbiter.scala 126:27]
  assign _GEN_20 = io_in_3_valid ? io_in_3_bits_way_en : _GEN_14; // @[Arbiter.scala 126:27]
  assign _GEN_21 = io_in_3_valid ? io_in_3_bits_idx : _GEN_15; // @[Arbiter.scala 126:27]
  assign _GEN_22 = io_in_3_valid ? io_in_3_bits_addr : _GEN_16; // @[Arbiter.scala 126:27]
  assign _GEN_23 = io_in_3_valid | io_in_4_valid; // @[Arbiter.scala 126:27]
  assign _GEN_25 = io_in_2_valid ? io_in_2_bits_data : _GEN_19; // @[Arbiter.scala 126:27]
  assign _GEN_26 = io_in_2_valid ? io_in_2_bits_way_en : _GEN_20; // @[Arbiter.scala 126:27]
  assign _GEN_27 = io_in_2_valid ? io_in_2_bits_idx : _GEN_21; // @[Arbiter.scala 126:27]
  assign _GEN_28 = io_in_2_valid ? io_in_2_bits_addr : _GEN_22; // @[Arbiter.scala 126:27]
  assign _GEN_29 = io_in_2_valid | _GEN_23; // @[Arbiter.scala 126:27]
  assign _T_210 = io_in_0_valid | io_in_2_valid; // @[Arbiter.scala 31:68]
  assign _T_211 = _T_210 | io_in_3_valid; // @[Arbiter.scala 31:68]
  assign _T_212 = _T_211 | io_in_4_valid; // @[Arbiter.scala 31:68]
  assign _T_213 = _T_212 | io_in_5_valid; // @[Arbiter.scala 31:68]
  assign _T_214 = _T_213 | io_in_6_valid; // @[Arbiter.scala 31:68]
  assign io_in_4_ready = ~_T_211 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_5_ready = ~_T_212 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_6_ready = ~_T_213 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_7_ready = ~_T_214 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = _T_214 | io_in_7_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_write = io_in_0_valid | _GEN_29; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_28; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_idx = io_in_0_valid ? io_in_0_bits_idx : _GEN_27; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_way_en = io_in_0_valid ? 4'hf : _GEN_26; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_data = io_in_0_valid ? io_in_0_bits_data : _GEN_25; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign Arbiter_covSum = 30'h0;
  assign io_covSum = Arbiter_covSum;
  assign metaAssert = 1'h0;
endmodule
module DCacheDataArray(
  input         clock,
  input         io_req_valid,
  input  [11:0] io_req_bits_addr,
  input         io_req_bits_write,
  input  [63:0] io_req_bits_wdata,
  input  [7:0]  io_req_bits_eccMask,
  input  [3:0]  io_req_bits_way_en,
  output [63:0] io_resp_0,
  output [63:0] io_resp_1,
  output [63:0] io_resp_2,
  output [63:0] io_resp_3,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [7:0] data_arrays_0_0 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_0;
  wire [7:0] data_arrays_0_0__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_0__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_0__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_0__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_0__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_0__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_0__T_211_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [8:0] data_arrays_0_0__T_211_addr_pipe_0;
  reg [31:0] _RAND_2;
  reg [7:0] data_arrays_0_1 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_3;
  wire [7:0] data_arrays_0_1__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_1__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_1__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_1__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_1__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_1__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_1__T_211_en_pipe_0;
  reg [31:0] _RAND_4;
  reg [8:0] data_arrays_0_1__T_211_addr_pipe_0;
  reg [31:0] _RAND_5;
  reg [7:0] data_arrays_0_2 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_6;
  wire [7:0] data_arrays_0_2__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_2__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_2__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_2__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_2__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_2__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_2__T_211_en_pipe_0;
  reg [31:0] _RAND_7;
  reg [8:0] data_arrays_0_2__T_211_addr_pipe_0;
  reg [31:0] _RAND_8;
  reg [7:0] data_arrays_0_3 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_9;
  wire [7:0] data_arrays_0_3__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_3__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_3__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_3__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_3__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_3__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_3__T_211_en_pipe_0;
  reg [31:0] _RAND_10;
  reg [8:0] data_arrays_0_3__T_211_addr_pipe_0;
  reg [31:0] _RAND_11;
  reg [7:0] data_arrays_0_4 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_12;
  wire [7:0] data_arrays_0_4__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_4__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_4__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_4__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_4__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_4__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_4__T_211_en_pipe_0;
  reg [31:0] _RAND_13;
  reg [8:0] data_arrays_0_4__T_211_addr_pipe_0;
  reg [31:0] _RAND_14;
  reg [7:0] data_arrays_0_5 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_15;
  wire [7:0] data_arrays_0_5__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_5__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_5__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_5__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_5__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_5__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_5__T_211_en_pipe_0;
  reg [31:0] _RAND_16;
  reg [8:0] data_arrays_0_5__T_211_addr_pipe_0;
  reg [31:0] _RAND_17;
  reg [7:0] data_arrays_0_6 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_18;
  wire [7:0] data_arrays_0_6__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_6__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_6__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_6__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_6__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_6__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_6__T_211_en_pipe_0;
  reg [31:0] _RAND_19;
  reg [8:0] data_arrays_0_6__T_211_addr_pipe_0;
  reg [31:0] _RAND_20;
  reg [7:0] data_arrays_0_7 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_21;
  wire [7:0] data_arrays_0_7__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_7__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_7__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_7__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_7__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_7__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_7__T_211_en_pipe_0;
  reg [31:0] _RAND_22;
  reg [8:0] data_arrays_0_7__T_211_addr_pipe_0;
  reg [31:0] _RAND_23;
  reg [7:0] data_arrays_0_8 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_24;
  wire [7:0] data_arrays_0_8__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_8__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_8__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_8__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_8__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_8__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_8__T_211_en_pipe_0;
  reg [31:0] _RAND_25;
  reg [8:0] data_arrays_0_8__T_211_addr_pipe_0;
  reg [31:0] _RAND_26;
  reg [7:0] data_arrays_0_9 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_27;
  wire [7:0] data_arrays_0_9__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_9__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_9__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_9__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_9__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_9__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_9__T_211_en_pipe_0;
  reg [31:0] _RAND_28;
  reg [8:0] data_arrays_0_9__T_211_addr_pipe_0;
  reg [31:0] _RAND_29;
  reg [7:0] data_arrays_0_10 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_30;
  wire [7:0] data_arrays_0_10__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_10__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_10__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_10__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_10__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_10__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_10__T_211_en_pipe_0;
  reg [31:0] _RAND_31;
  reg [8:0] data_arrays_0_10__T_211_addr_pipe_0;
  reg [31:0] _RAND_32;
  reg [7:0] data_arrays_0_11 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_33;
  wire [7:0] data_arrays_0_11__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_11__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_11__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_11__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_11__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_11__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_11__T_211_en_pipe_0;
  reg [31:0] _RAND_34;
  reg [8:0] data_arrays_0_11__T_211_addr_pipe_0;
  reg [31:0] _RAND_35;
  reg [7:0] data_arrays_0_12 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_36;
  wire [7:0] data_arrays_0_12__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_12__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_12__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_12__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_12__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_12__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_12__T_211_en_pipe_0;
  reg [31:0] _RAND_37;
  reg [8:0] data_arrays_0_12__T_211_addr_pipe_0;
  reg [31:0] _RAND_38;
  reg [7:0] data_arrays_0_13 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_39;
  wire [7:0] data_arrays_0_13__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_13__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_13__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_13__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_13__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_13__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_13__T_211_en_pipe_0;
  reg [31:0] _RAND_40;
  reg [8:0] data_arrays_0_13__T_211_addr_pipe_0;
  reg [31:0] _RAND_41;
  reg [7:0] data_arrays_0_14 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_42;
  wire [7:0] data_arrays_0_14__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_14__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_14__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_14__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_14__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_14__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_14__T_211_en_pipe_0;
  reg [31:0] _RAND_43;
  reg [8:0] data_arrays_0_14__T_211_addr_pipe_0;
  reg [31:0] _RAND_44;
  reg [7:0] data_arrays_0_15 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_45;
  wire [7:0] data_arrays_0_15__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_15__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_15__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_15__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_15__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_15__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_15__T_211_en_pipe_0;
  reg [31:0] _RAND_46;
  reg [8:0] data_arrays_0_15__T_211_addr_pipe_0;
  reg [31:0] _RAND_47;
  reg [7:0] data_arrays_0_16 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_48;
  wire [7:0] data_arrays_0_16__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_16__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_16__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_16__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_16__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_16__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_16__T_211_en_pipe_0;
  reg [31:0] _RAND_49;
  reg [8:0] data_arrays_0_16__T_211_addr_pipe_0;
  reg [31:0] _RAND_50;
  reg [7:0] data_arrays_0_17 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_51;
  wire [7:0] data_arrays_0_17__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_17__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_17__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_17__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_17__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_17__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_17__T_211_en_pipe_0;
  reg [31:0] _RAND_52;
  reg [8:0] data_arrays_0_17__T_211_addr_pipe_0;
  reg [31:0] _RAND_53;
  reg [7:0] data_arrays_0_18 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_54;
  wire [7:0] data_arrays_0_18__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_18__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_18__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_18__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_18__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_18__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_18__T_211_en_pipe_0;
  reg [31:0] _RAND_55;
  reg [8:0] data_arrays_0_18__T_211_addr_pipe_0;
  reg [31:0] _RAND_56;
  reg [7:0] data_arrays_0_19 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_57;
  wire [7:0] data_arrays_0_19__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_19__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_19__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_19__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_19__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_19__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_19__T_211_en_pipe_0;
  reg [31:0] _RAND_58;
  reg [8:0] data_arrays_0_19__T_211_addr_pipe_0;
  reg [31:0] _RAND_59;
  reg [7:0] data_arrays_0_20 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_60;
  wire [7:0] data_arrays_0_20__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_20__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_20__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_20__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_20__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_20__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_20__T_211_en_pipe_0;
  reg [31:0] _RAND_61;
  reg [8:0] data_arrays_0_20__T_211_addr_pipe_0;
  reg [31:0] _RAND_62;
  reg [7:0] data_arrays_0_21 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_63;
  wire [7:0] data_arrays_0_21__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_21__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_21__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_21__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_21__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_21__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_21__T_211_en_pipe_0;
  reg [31:0] _RAND_64;
  reg [8:0] data_arrays_0_21__T_211_addr_pipe_0;
  reg [31:0] _RAND_65;
  reg [7:0] data_arrays_0_22 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_66;
  wire [7:0] data_arrays_0_22__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_22__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_22__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_22__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_22__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_22__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_22__T_211_en_pipe_0;
  reg [31:0] _RAND_67;
  reg [8:0] data_arrays_0_22__T_211_addr_pipe_0;
  reg [31:0] _RAND_68;
  reg [7:0] data_arrays_0_23 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_69;
  wire [7:0] data_arrays_0_23__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_23__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_23__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_23__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_23__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_23__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_23__T_211_en_pipe_0;
  reg [31:0] _RAND_70;
  reg [8:0] data_arrays_0_23__T_211_addr_pipe_0;
  reg [31:0] _RAND_71;
  reg [7:0] data_arrays_0_24 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_72;
  wire [7:0] data_arrays_0_24__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_24__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_24__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_24__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_24__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_24__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_24__T_211_en_pipe_0;
  reg [31:0] _RAND_73;
  reg [8:0] data_arrays_0_24__T_211_addr_pipe_0;
  reg [31:0] _RAND_74;
  reg [7:0] data_arrays_0_25 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_75;
  wire [7:0] data_arrays_0_25__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_25__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_25__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_25__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_25__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_25__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_25__T_211_en_pipe_0;
  reg [31:0] _RAND_76;
  reg [8:0] data_arrays_0_25__T_211_addr_pipe_0;
  reg [31:0] _RAND_77;
  reg [7:0] data_arrays_0_26 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_78;
  wire [7:0] data_arrays_0_26__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_26__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_26__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_26__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_26__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_26__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_26__T_211_en_pipe_0;
  reg [31:0] _RAND_79;
  reg [8:0] data_arrays_0_26__T_211_addr_pipe_0;
  reg [31:0] _RAND_80;
  reg [7:0] data_arrays_0_27 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_81;
  wire [7:0] data_arrays_0_27__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_27__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_27__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_27__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_27__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_27__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_27__T_211_en_pipe_0;
  reg [31:0] _RAND_82;
  reg [8:0] data_arrays_0_27__T_211_addr_pipe_0;
  reg [31:0] _RAND_83;
  reg [7:0] data_arrays_0_28 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_84;
  wire [7:0] data_arrays_0_28__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_28__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_28__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_28__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_28__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_28__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_28__T_211_en_pipe_0;
  reg [31:0] _RAND_85;
  reg [8:0] data_arrays_0_28__T_211_addr_pipe_0;
  reg [31:0] _RAND_86;
  reg [7:0] data_arrays_0_29 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_87;
  wire [7:0] data_arrays_0_29__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_29__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_29__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_29__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_29__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_29__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_29__T_211_en_pipe_0;
  reg [31:0] _RAND_88;
  reg [8:0] data_arrays_0_29__T_211_addr_pipe_0;
  reg [31:0] _RAND_89;
  reg [7:0] data_arrays_0_30 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_90;
  wire [7:0] data_arrays_0_30__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_30__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_30__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_30__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_30__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_30__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_30__T_211_en_pipe_0;
  reg [31:0] _RAND_91;
  reg [8:0] data_arrays_0_30__T_211_addr_pipe_0;
  reg [31:0] _RAND_92;
  reg [7:0] data_arrays_0_31 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_93;
  wire [7:0] data_arrays_0_31__T_211_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_31__T_211_addr; // @[DescribedSRAM.scala 23:21]
  wire [7:0] data_arrays_0_31__T_137_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_31__T_137_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_31__T_137_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_31__T_137_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_31__T_211_en_pipe_0;
  reg [31:0] _RAND_94;
  reg [8:0] data_arrays_0_31__T_211_addr_pipe_0;
  reg [31:0] _RAND_95;
  wire  eccMask_0; // @[DCache.scala 41:79]
  wire  eccMask_1; // @[DCache.scala 41:79]
  wire  eccMask_2; // @[DCache.scala 41:79]
  wire  eccMask_3; // @[DCache.scala 41:79]
  wire  eccMask_4; // @[DCache.scala 41:79]
  wire  eccMask_5; // @[DCache.scala 41:79]
  wire  eccMask_6; // @[DCache.scala 41:79]
  wire  eccMask_7; // @[DCache.scala 41:79]
  wire [31:0] _T_281; // @[Cat.scala 30:58]
  wire [31:0] _T_284; // @[Cat.scala 30:58]
  wire [31:0] _T_287; // @[Cat.scala 30:58]
  wire [31:0] _T_290; // @[Cat.scala 30:58]
  wire [31:0] _T_293; // @[Cat.scala 30:58]
  wire [31:0] _T_296; // @[Cat.scala 30:58]
  wire [31:0] _T_299; // @[Cat.scala 30:58]
  wire [31:0] _T_302; // @[Cat.scala 30:58]
  wire [29:0] DCacheDataArray_covSum;
  assign data_arrays_0_0__T_211_addr = data_arrays_0_0__T_211_addr_pipe_0;
  assign data_arrays_0_0__T_211_data = data_arrays_0_0[data_arrays_0_0__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_0__T_137_data = io_req_bits_wdata[7:0];
  assign data_arrays_0_0__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_0__T_137_mask = eccMask_0 & io_req_bits_way_en[0];
  assign data_arrays_0_0__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_1__T_211_addr = data_arrays_0_1__T_211_addr_pipe_0;
  assign data_arrays_0_1__T_211_data = data_arrays_0_1[data_arrays_0_1__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_1__T_137_data = io_req_bits_wdata[15:8];
  assign data_arrays_0_1__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_1__T_137_mask = eccMask_1 & io_req_bits_way_en[0];
  assign data_arrays_0_1__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_2__T_211_addr = data_arrays_0_2__T_211_addr_pipe_0;
  assign data_arrays_0_2__T_211_data = data_arrays_0_2[data_arrays_0_2__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_2__T_137_data = io_req_bits_wdata[23:16];
  assign data_arrays_0_2__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_2__T_137_mask = eccMask_2 & io_req_bits_way_en[0];
  assign data_arrays_0_2__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_3__T_211_addr = data_arrays_0_3__T_211_addr_pipe_0;
  assign data_arrays_0_3__T_211_data = data_arrays_0_3[data_arrays_0_3__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_3__T_137_data = io_req_bits_wdata[31:24];
  assign data_arrays_0_3__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_3__T_137_mask = eccMask_3 & io_req_bits_way_en[0];
  assign data_arrays_0_3__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_4__T_211_addr = data_arrays_0_4__T_211_addr_pipe_0;
  assign data_arrays_0_4__T_211_data = data_arrays_0_4[data_arrays_0_4__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_4__T_137_data = io_req_bits_wdata[39:32];
  assign data_arrays_0_4__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_4__T_137_mask = eccMask_4 & io_req_bits_way_en[0];
  assign data_arrays_0_4__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_5__T_211_addr = data_arrays_0_5__T_211_addr_pipe_0;
  assign data_arrays_0_5__T_211_data = data_arrays_0_5[data_arrays_0_5__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_5__T_137_data = io_req_bits_wdata[47:40];
  assign data_arrays_0_5__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_5__T_137_mask = eccMask_5 & io_req_bits_way_en[0];
  assign data_arrays_0_5__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_6__T_211_addr = data_arrays_0_6__T_211_addr_pipe_0;
  assign data_arrays_0_6__T_211_data = data_arrays_0_6[data_arrays_0_6__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_6__T_137_data = io_req_bits_wdata[55:48];
  assign data_arrays_0_6__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_6__T_137_mask = eccMask_6 & io_req_bits_way_en[0];
  assign data_arrays_0_6__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_7__T_211_addr = data_arrays_0_7__T_211_addr_pipe_0;
  assign data_arrays_0_7__T_211_data = data_arrays_0_7[data_arrays_0_7__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_7__T_137_data = io_req_bits_wdata[63:56];
  assign data_arrays_0_7__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_7__T_137_mask = eccMask_7 & io_req_bits_way_en[0];
  assign data_arrays_0_7__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_8__T_211_addr = data_arrays_0_8__T_211_addr_pipe_0;
  assign data_arrays_0_8__T_211_data = data_arrays_0_8[data_arrays_0_8__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_8__T_137_data = io_req_bits_wdata[7:0];
  assign data_arrays_0_8__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_8__T_137_mask = eccMask_0 & io_req_bits_way_en[1];
  assign data_arrays_0_8__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_9__T_211_addr = data_arrays_0_9__T_211_addr_pipe_0;
  assign data_arrays_0_9__T_211_data = data_arrays_0_9[data_arrays_0_9__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_9__T_137_data = io_req_bits_wdata[15:8];
  assign data_arrays_0_9__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_9__T_137_mask = eccMask_1 & io_req_bits_way_en[1];
  assign data_arrays_0_9__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_10__T_211_addr = data_arrays_0_10__T_211_addr_pipe_0;
  assign data_arrays_0_10__T_211_data = data_arrays_0_10[data_arrays_0_10__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_10__T_137_data = io_req_bits_wdata[23:16];
  assign data_arrays_0_10__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_10__T_137_mask = eccMask_2 & io_req_bits_way_en[1];
  assign data_arrays_0_10__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_11__T_211_addr = data_arrays_0_11__T_211_addr_pipe_0;
  assign data_arrays_0_11__T_211_data = data_arrays_0_11[data_arrays_0_11__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_11__T_137_data = io_req_bits_wdata[31:24];
  assign data_arrays_0_11__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_11__T_137_mask = eccMask_3 & io_req_bits_way_en[1];
  assign data_arrays_0_11__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_12__T_211_addr = data_arrays_0_12__T_211_addr_pipe_0;
  assign data_arrays_0_12__T_211_data = data_arrays_0_12[data_arrays_0_12__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_12__T_137_data = io_req_bits_wdata[39:32];
  assign data_arrays_0_12__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_12__T_137_mask = eccMask_4 & io_req_bits_way_en[1];
  assign data_arrays_0_12__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_13__T_211_addr = data_arrays_0_13__T_211_addr_pipe_0;
  assign data_arrays_0_13__T_211_data = data_arrays_0_13[data_arrays_0_13__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_13__T_137_data = io_req_bits_wdata[47:40];
  assign data_arrays_0_13__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_13__T_137_mask = eccMask_5 & io_req_bits_way_en[1];
  assign data_arrays_0_13__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_14__T_211_addr = data_arrays_0_14__T_211_addr_pipe_0;
  assign data_arrays_0_14__T_211_data = data_arrays_0_14[data_arrays_0_14__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_14__T_137_data = io_req_bits_wdata[55:48];
  assign data_arrays_0_14__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_14__T_137_mask = eccMask_6 & io_req_bits_way_en[1];
  assign data_arrays_0_14__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_15__T_211_addr = data_arrays_0_15__T_211_addr_pipe_0;
  assign data_arrays_0_15__T_211_data = data_arrays_0_15[data_arrays_0_15__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_15__T_137_data = io_req_bits_wdata[63:56];
  assign data_arrays_0_15__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_15__T_137_mask = eccMask_7 & io_req_bits_way_en[1];
  assign data_arrays_0_15__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_16__T_211_addr = data_arrays_0_16__T_211_addr_pipe_0;
  assign data_arrays_0_16__T_211_data = data_arrays_0_16[data_arrays_0_16__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_16__T_137_data = io_req_bits_wdata[7:0];
  assign data_arrays_0_16__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_16__T_137_mask = eccMask_0 & io_req_bits_way_en[2];
  assign data_arrays_0_16__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_17__T_211_addr = data_arrays_0_17__T_211_addr_pipe_0;
  assign data_arrays_0_17__T_211_data = data_arrays_0_17[data_arrays_0_17__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_17__T_137_data = io_req_bits_wdata[15:8];
  assign data_arrays_0_17__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_17__T_137_mask = eccMask_1 & io_req_bits_way_en[2];
  assign data_arrays_0_17__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_18__T_211_addr = data_arrays_0_18__T_211_addr_pipe_0;
  assign data_arrays_0_18__T_211_data = data_arrays_0_18[data_arrays_0_18__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_18__T_137_data = io_req_bits_wdata[23:16];
  assign data_arrays_0_18__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_18__T_137_mask = eccMask_2 & io_req_bits_way_en[2];
  assign data_arrays_0_18__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_19__T_211_addr = data_arrays_0_19__T_211_addr_pipe_0;
  assign data_arrays_0_19__T_211_data = data_arrays_0_19[data_arrays_0_19__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_19__T_137_data = io_req_bits_wdata[31:24];
  assign data_arrays_0_19__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_19__T_137_mask = eccMask_3 & io_req_bits_way_en[2];
  assign data_arrays_0_19__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_20__T_211_addr = data_arrays_0_20__T_211_addr_pipe_0;
  assign data_arrays_0_20__T_211_data = data_arrays_0_20[data_arrays_0_20__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_20__T_137_data = io_req_bits_wdata[39:32];
  assign data_arrays_0_20__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_20__T_137_mask = eccMask_4 & io_req_bits_way_en[2];
  assign data_arrays_0_20__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_21__T_211_addr = data_arrays_0_21__T_211_addr_pipe_0;
  assign data_arrays_0_21__T_211_data = data_arrays_0_21[data_arrays_0_21__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_21__T_137_data = io_req_bits_wdata[47:40];
  assign data_arrays_0_21__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_21__T_137_mask = eccMask_5 & io_req_bits_way_en[2];
  assign data_arrays_0_21__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_22__T_211_addr = data_arrays_0_22__T_211_addr_pipe_0;
  assign data_arrays_0_22__T_211_data = data_arrays_0_22[data_arrays_0_22__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_22__T_137_data = io_req_bits_wdata[55:48];
  assign data_arrays_0_22__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_22__T_137_mask = eccMask_6 & io_req_bits_way_en[2];
  assign data_arrays_0_22__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_23__T_211_addr = data_arrays_0_23__T_211_addr_pipe_0;
  assign data_arrays_0_23__T_211_data = data_arrays_0_23[data_arrays_0_23__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_23__T_137_data = io_req_bits_wdata[63:56];
  assign data_arrays_0_23__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_23__T_137_mask = eccMask_7 & io_req_bits_way_en[2];
  assign data_arrays_0_23__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_24__T_211_addr = data_arrays_0_24__T_211_addr_pipe_0;
  assign data_arrays_0_24__T_211_data = data_arrays_0_24[data_arrays_0_24__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_24__T_137_data = io_req_bits_wdata[7:0];
  assign data_arrays_0_24__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_24__T_137_mask = eccMask_0 & io_req_bits_way_en[3];
  assign data_arrays_0_24__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_25__T_211_addr = data_arrays_0_25__T_211_addr_pipe_0;
  assign data_arrays_0_25__T_211_data = data_arrays_0_25[data_arrays_0_25__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_25__T_137_data = io_req_bits_wdata[15:8];
  assign data_arrays_0_25__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_25__T_137_mask = eccMask_1 & io_req_bits_way_en[3];
  assign data_arrays_0_25__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_26__T_211_addr = data_arrays_0_26__T_211_addr_pipe_0;
  assign data_arrays_0_26__T_211_data = data_arrays_0_26[data_arrays_0_26__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_26__T_137_data = io_req_bits_wdata[23:16];
  assign data_arrays_0_26__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_26__T_137_mask = eccMask_2 & io_req_bits_way_en[3];
  assign data_arrays_0_26__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_27__T_211_addr = data_arrays_0_27__T_211_addr_pipe_0;
  assign data_arrays_0_27__T_211_data = data_arrays_0_27[data_arrays_0_27__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_27__T_137_data = io_req_bits_wdata[31:24];
  assign data_arrays_0_27__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_27__T_137_mask = eccMask_3 & io_req_bits_way_en[3];
  assign data_arrays_0_27__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_28__T_211_addr = data_arrays_0_28__T_211_addr_pipe_0;
  assign data_arrays_0_28__T_211_data = data_arrays_0_28[data_arrays_0_28__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_28__T_137_data = io_req_bits_wdata[39:32];
  assign data_arrays_0_28__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_28__T_137_mask = eccMask_4 & io_req_bits_way_en[3];
  assign data_arrays_0_28__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_29__T_211_addr = data_arrays_0_29__T_211_addr_pipe_0;
  assign data_arrays_0_29__T_211_data = data_arrays_0_29[data_arrays_0_29__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_29__T_137_data = io_req_bits_wdata[47:40];
  assign data_arrays_0_29__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_29__T_137_mask = eccMask_5 & io_req_bits_way_en[3];
  assign data_arrays_0_29__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_30__T_211_addr = data_arrays_0_30__T_211_addr_pipe_0;
  assign data_arrays_0_30__T_211_data = data_arrays_0_30[data_arrays_0_30__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_30__T_137_data = io_req_bits_wdata[55:48];
  assign data_arrays_0_30__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_30__T_137_mask = eccMask_6 & io_req_bits_way_en[3];
  assign data_arrays_0_30__T_137_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_31__T_211_addr = data_arrays_0_31__T_211_addr_pipe_0;
  assign data_arrays_0_31__T_211_data = data_arrays_0_31[data_arrays_0_31__T_211_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_31__T_137_data = io_req_bits_wdata[63:56];
  assign data_arrays_0_31__T_137_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_31__T_137_mask = eccMask_7 & io_req_bits_way_en[3];
  assign data_arrays_0_31__T_137_en = io_req_valid & io_req_bits_write;
  assign eccMask_0 = io_req_bits_eccMask[0]; // @[DCache.scala 41:79]
  assign eccMask_1 = io_req_bits_eccMask[1]; // @[DCache.scala 41:79]
  assign eccMask_2 = io_req_bits_eccMask[2]; // @[DCache.scala 41:79]
  assign eccMask_3 = io_req_bits_eccMask[3]; // @[DCache.scala 41:79]
  assign eccMask_4 = io_req_bits_eccMask[4]; // @[DCache.scala 41:79]
  assign eccMask_5 = io_req_bits_eccMask[5]; // @[DCache.scala 41:79]
  assign eccMask_6 = io_req_bits_eccMask[6]; // @[DCache.scala 41:79]
  assign eccMask_7 = io_req_bits_eccMask[7]; // @[DCache.scala 41:79]
  assign _T_281 = {data_arrays_0_3__T_211_data,data_arrays_0_2__T_211_data,data_arrays_0_1__T_211_data,data_arrays_0_0__T_211_data}; // @[Cat.scala 30:58]
  assign _T_284 = {data_arrays_0_7__T_211_data,data_arrays_0_6__T_211_data,data_arrays_0_5__T_211_data,data_arrays_0_4__T_211_data}; // @[Cat.scala 30:58]
  assign _T_287 = {data_arrays_0_11__T_211_data,data_arrays_0_10__T_211_data,data_arrays_0_9__T_211_data,data_arrays_0_8__T_211_data}; // @[Cat.scala 30:58]
  assign _T_290 = {data_arrays_0_15__T_211_data,data_arrays_0_14__T_211_data,data_arrays_0_13__T_211_data,data_arrays_0_12__T_211_data}; // @[Cat.scala 30:58]
  assign _T_293 = {data_arrays_0_19__T_211_data,data_arrays_0_18__T_211_data,data_arrays_0_17__T_211_data,data_arrays_0_16__T_211_data}; // @[Cat.scala 30:58]
  assign _T_296 = {data_arrays_0_23__T_211_data,data_arrays_0_22__T_211_data,data_arrays_0_21__T_211_data,data_arrays_0_20__T_211_data}; // @[Cat.scala 30:58]
  assign _T_299 = {data_arrays_0_27__T_211_data,data_arrays_0_26__T_211_data,data_arrays_0_25__T_211_data,data_arrays_0_24__T_211_data}; // @[Cat.scala 30:58]
  assign _T_302 = {data_arrays_0_31__T_211_data,data_arrays_0_30__T_211_data,data_arrays_0_29__T_211_data,data_arrays_0_28__T_211_data}; // @[Cat.scala 30:58]
  assign io_resp_0 = {_T_284,_T_281}; // @[DCache.scala 64:69]
  assign io_resp_1 = {_T_290,_T_287}; // @[DCache.scala 64:69]
  assign io_resp_2 = {_T_296,_T_293}; // @[DCache.scala 64:69]
  assign io_resp_3 = {_T_302,_T_299}; // @[DCache.scala 64:69]
  assign DCacheDataArray_covSum = 30'h0;
  assign io_covSum = DCacheDataArray_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_0[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  data_arrays_0_0__T_211_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  data_arrays_0_0__T_211_addr_pipe_0 = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_1[initvar] = _RAND_3[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  data_arrays_0_1__T_211_en_pipe_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  data_arrays_0_1__T_211_addr_pipe_0 = _RAND_5[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_2[initvar] = _RAND_6[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  data_arrays_0_2__T_211_en_pipe_0 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  data_arrays_0_2__T_211_addr_pipe_0 = _RAND_8[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_3[initvar] = _RAND_9[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_arrays_0_3__T_211_en_pipe_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  data_arrays_0_3__T_211_addr_pipe_0 = _RAND_11[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_4[initvar] = _RAND_12[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  data_arrays_0_4__T_211_en_pipe_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  data_arrays_0_4__T_211_addr_pipe_0 = _RAND_14[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_5[initvar] = _RAND_15[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  data_arrays_0_5__T_211_en_pipe_0 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  data_arrays_0_5__T_211_addr_pipe_0 = _RAND_17[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_6[initvar] = _RAND_18[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  data_arrays_0_6__T_211_en_pipe_0 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  data_arrays_0_6__T_211_addr_pipe_0 = _RAND_20[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_7[initvar] = _RAND_21[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  data_arrays_0_7__T_211_en_pipe_0 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  data_arrays_0_7__T_211_addr_pipe_0 = _RAND_23[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_8[initvar] = _RAND_24[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  data_arrays_0_8__T_211_en_pipe_0 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  data_arrays_0_8__T_211_addr_pipe_0 = _RAND_26[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_9[initvar] = _RAND_27[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  data_arrays_0_9__T_211_en_pipe_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  data_arrays_0_9__T_211_addr_pipe_0 = _RAND_29[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_10[initvar] = _RAND_30[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  data_arrays_0_10__T_211_en_pipe_0 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  data_arrays_0_10__T_211_addr_pipe_0 = _RAND_32[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_11[initvar] = _RAND_33[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  data_arrays_0_11__T_211_en_pipe_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  data_arrays_0_11__T_211_addr_pipe_0 = _RAND_35[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_12[initvar] = _RAND_36[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  data_arrays_0_12__T_211_en_pipe_0 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  data_arrays_0_12__T_211_addr_pipe_0 = _RAND_38[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_13[initvar] = _RAND_39[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  data_arrays_0_13__T_211_en_pipe_0 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  data_arrays_0_13__T_211_addr_pipe_0 = _RAND_41[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_14[initvar] = _RAND_42[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  data_arrays_0_14__T_211_en_pipe_0 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  data_arrays_0_14__T_211_addr_pipe_0 = _RAND_44[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_15[initvar] = _RAND_45[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  data_arrays_0_15__T_211_en_pipe_0 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  data_arrays_0_15__T_211_addr_pipe_0 = _RAND_47[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_16[initvar] = _RAND_48[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  data_arrays_0_16__T_211_en_pipe_0 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  data_arrays_0_16__T_211_addr_pipe_0 = _RAND_50[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_17[initvar] = _RAND_51[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  data_arrays_0_17__T_211_en_pipe_0 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  data_arrays_0_17__T_211_addr_pipe_0 = _RAND_53[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_18[initvar] = _RAND_54[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  data_arrays_0_18__T_211_en_pipe_0 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  data_arrays_0_18__T_211_addr_pipe_0 = _RAND_56[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_19[initvar] = _RAND_57[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  data_arrays_0_19__T_211_en_pipe_0 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  data_arrays_0_19__T_211_addr_pipe_0 = _RAND_59[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_20[initvar] = _RAND_60[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  data_arrays_0_20__T_211_en_pipe_0 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  data_arrays_0_20__T_211_addr_pipe_0 = _RAND_62[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_21[initvar] = _RAND_63[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  data_arrays_0_21__T_211_en_pipe_0 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  data_arrays_0_21__T_211_addr_pipe_0 = _RAND_65[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_22[initvar] = _RAND_66[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  data_arrays_0_22__T_211_en_pipe_0 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  data_arrays_0_22__T_211_addr_pipe_0 = _RAND_68[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_23[initvar] = _RAND_69[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  data_arrays_0_23__T_211_en_pipe_0 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  data_arrays_0_23__T_211_addr_pipe_0 = _RAND_71[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_24[initvar] = _RAND_72[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  data_arrays_0_24__T_211_en_pipe_0 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  data_arrays_0_24__T_211_addr_pipe_0 = _RAND_74[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_25[initvar] = _RAND_75[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  data_arrays_0_25__T_211_en_pipe_0 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  data_arrays_0_25__T_211_addr_pipe_0 = _RAND_77[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_26[initvar] = _RAND_78[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  data_arrays_0_26__T_211_en_pipe_0 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  data_arrays_0_26__T_211_addr_pipe_0 = _RAND_80[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_27[initvar] = _RAND_81[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  data_arrays_0_27__T_211_en_pipe_0 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  data_arrays_0_27__T_211_addr_pipe_0 = _RAND_83[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_28[initvar] = _RAND_84[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  data_arrays_0_28__T_211_en_pipe_0 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  data_arrays_0_28__T_211_addr_pipe_0 = _RAND_86[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_29[initvar] = _RAND_87[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  data_arrays_0_29__T_211_en_pipe_0 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  data_arrays_0_29__T_211_addr_pipe_0 = _RAND_89[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_30[initvar] = _RAND_90[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  data_arrays_0_30__T_211_en_pipe_0 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  data_arrays_0_30__T_211_addr_pipe_0 = _RAND_92[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_31[initvar] = _RAND_93[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  data_arrays_0_31__T_211_en_pipe_0 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  data_arrays_0_31__T_211_addr_pipe_0 = _RAND_95[8:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(data_arrays_0_0__T_137_en & data_arrays_0_0__T_137_mask) begin
      data_arrays_0_0[data_arrays_0_0__T_137_addr] <= data_arrays_0_0__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_0__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_0__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_0__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_0__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_1__T_137_en & data_arrays_0_1__T_137_mask) begin
      data_arrays_0_1[data_arrays_0_1__T_137_addr] <= data_arrays_0_1__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_1__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_1__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_1__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_1__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_2__T_137_en & data_arrays_0_2__T_137_mask) begin
      data_arrays_0_2[data_arrays_0_2__T_137_addr] <= data_arrays_0_2__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_2__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_2__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_2__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_2__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_3__T_137_en & data_arrays_0_3__T_137_mask) begin
      data_arrays_0_3[data_arrays_0_3__T_137_addr] <= data_arrays_0_3__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_3__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_3__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_3__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_3__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_4__T_137_en & data_arrays_0_4__T_137_mask) begin
      data_arrays_0_4[data_arrays_0_4__T_137_addr] <= data_arrays_0_4__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_4__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_4__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_4__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_4__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_5__T_137_en & data_arrays_0_5__T_137_mask) begin
      data_arrays_0_5[data_arrays_0_5__T_137_addr] <= data_arrays_0_5__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_5__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_5__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_5__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_5__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_6__T_137_en & data_arrays_0_6__T_137_mask) begin
      data_arrays_0_6[data_arrays_0_6__T_137_addr] <= data_arrays_0_6__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_6__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_6__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_6__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_6__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_7__T_137_en & data_arrays_0_7__T_137_mask) begin
      data_arrays_0_7[data_arrays_0_7__T_137_addr] <= data_arrays_0_7__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_7__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_7__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_7__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_7__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_8__T_137_en & data_arrays_0_8__T_137_mask) begin
      data_arrays_0_8[data_arrays_0_8__T_137_addr] <= data_arrays_0_8__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_8__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_8__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_8__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_8__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_9__T_137_en & data_arrays_0_9__T_137_mask) begin
      data_arrays_0_9[data_arrays_0_9__T_137_addr] <= data_arrays_0_9__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_9__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_9__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_9__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_9__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_10__T_137_en & data_arrays_0_10__T_137_mask) begin
      data_arrays_0_10[data_arrays_0_10__T_137_addr] <= data_arrays_0_10__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_10__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_10__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_10__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_10__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_11__T_137_en & data_arrays_0_11__T_137_mask) begin
      data_arrays_0_11[data_arrays_0_11__T_137_addr] <= data_arrays_0_11__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_11__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_11__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_11__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_11__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_12__T_137_en & data_arrays_0_12__T_137_mask) begin
      data_arrays_0_12[data_arrays_0_12__T_137_addr] <= data_arrays_0_12__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_12__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_12__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_12__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_12__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_13__T_137_en & data_arrays_0_13__T_137_mask) begin
      data_arrays_0_13[data_arrays_0_13__T_137_addr] <= data_arrays_0_13__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_13__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_13__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_13__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_13__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_14__T_137_en & data_arrays_0_14__T_137_mask) begin
      data_arrays_0_14[data_arrays_0_14__T_137_addr] <= data_arrays_0_14__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_14__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_14__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_14__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_14__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_15__T_137_en & data_arrays_0_15__T_137_mask) begin
      data_arrays_0_15[data_arrays_0_15__T_137_addr] <= data_arrays_0_15__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_15__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_15__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_15__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_15__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_16__T_137_en & data_arrays_0_16__T_137_mask) begin
      data_arrays_0_16[data_arrays_0_16__T_137_addr] <= data_arrays_0_16__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_16__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_16__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_16__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_16__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_17__T_137_en & data_arrays_0_17__T_137_mask) begin
      data_arrays_0_17[data_arrays_0_17__T_137_addr] <= data_arrays_0_17__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_17__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_17__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_17__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_17__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_18__T_137_en & data_arrays_0_18__T_137_mask) begin
      data_arrays_0_18[data_arrays_0_18__T_137_addr] <= data_arrays_0_18__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_18__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_18__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_18__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_18__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_19__T_137_en & data_arrays_0_19__T_137_mask) begin
      data_arrays_0_19[data_arrays_0_19__T_137_addr] <= data_arrays_0_19__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_19__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_19__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_19__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_19__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_20__T_137_en & data_arrays_0_20__T_137_mask) begin
      data_arrays_0_20[data_arrays_0_20__T_137_addr] <= data_arrays_0_20__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_20__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_20__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_20__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_20__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_21__T_137_en & data_arrays_0_21__T_137_mask) begin
      data_arrays_0_21[data_arrays_0_21__T_137_addr] <= data_arrays_0_21__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_21__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_21__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_21__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_21__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_22__T_137_en & data_arrays_0_22__T_137_mask) begin
      data_arrays_0_22[data_arrays_0_22__T_137_addr] <= data_arrays_0_22__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_22__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_22__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_22__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_22__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_23__T_137_en & data_arrays_0_23__T_137_mask) begin
      data_arrays_0_23[data_arrays_0_23__T_137_addr] <= data_arrays_0_23__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_23__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_23__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_23__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_23__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_24__T_137_en & data_arrays_0_24__T_137_mask) begin
      data_arrays_0_24[data_arrays_0_24__T_137_addr] <= data_arrays_0_24__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_24__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_24__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_24__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_24__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_25__T_137_en & data_arrays_0_25__T_137_mask) begin
      data_arrays_0_25[data_arrays_0_25__T_137_addr] <= data_arrays_0_25__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_25__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_25__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_25__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_25__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_26__T_137_en & data_arrays_0_26__T_137_mask) begin
      data_arrays_0_26[data_arrays_0_26__T_137_addr] <= data_arrays_0_26__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_26__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_26__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_26__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_26__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_27__T_137_en & data_arrays_0_27__T_137_mask) begin
      data_arrays_0_27[data_arrays_0_27__T_137_addr] <= data_arrays_0_27__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_27__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_27__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_27__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_27__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_28__T_137_en & data_arrays_0_28__T_137_mask) begin
      data_arrays_0_28[data_arrays_0_28__T_137_addr] <= data_arrays_0_28__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_28__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_28__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_28__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_28__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_29__T_137_en & data_arrays_0_29__T_137_mask) begin
      data_arrays_0_29[data_arrays_0_29__T_137_addr] <= data_arrays_0_29__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_29__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_29__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_29__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_29__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_30__T_137_en & data_arrays_0_30__T_137_mask) begin
      data_arrays_0_30[data_arrays_0_30__T_137_addr] <= data_arrays_0_30__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_30__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_30__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_30__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_30__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_31__T_137_en & data_arrays_0_31__T_137_mask) begin
      data_arrays_0_31[data_arrays_0_31__T_137_addr] <= data_arrays_0_31__T_137_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_31__T_211_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_31__T_211_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_31__T_211_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_31__T_211_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
  end
endmodule
module Arbiter_1(
  input         io_in_0_valid,
  input  [11:0] io_in_0_bits_addr,
  input         io_in_0_bits_write,
  input  [63:0] io_in_0_bits_wdata,
  input  [7:0]  io_in_0_bits_eccMask,
  input  [3:0]  io_in_0_bits_way_en,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [11:0] io_in_1_bits_addr,
  input         io_in_1_bits_write,
  input  [63:0] io_in_1_bits_wdata,
  input  [7:0]  io_in_1_bits_eccMask,
  input  [3:0]  io_in_1_bits_way_en,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [11:0] io_in_2_bits_addr,
  input  [63:0] io_in_2_bits_wdata,
  input  [7:0]  io_in_2_bits_eccMask,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input  [11:0] io_in_3_bits_addr,
  input  [63:0] io_in_3_bits_wdata,
  input  [7:0]  io_in_3_bits_eccMask,
  output        io_out_valid,
  output [11:0] io_out_bits_addr,
  output        io_out_bits_write,
  output [63:0] io_out_bits_wdata,
  output [7:0]  io_out_bits_eccMask,
  output [3:0]  io_out_bits_way_en,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [7:0] _GEN_2; // @[Arbiter.scala 126:27]
  wire [63:0] _GEN_5; // @[Arbiter.scala 126:27]
  wire [11:0] _GEN_7; // @[Arbiter.scala 126:27]
  wire [3:0] _GEN_9; // @[Arbiter.scala 126:27]
  wire [7:0] _GEN_10; // @[Arbiter.scala 126:27]
  wire [63:0] _GEN_13; // @[Arbiter.scala 126:27]
  wire  _GEN_14; // @[Arbiter.scala 126:27]
  wire [11:0] _GEN_15; // @[Arbiter.scala 126:27]
  wire  _T_94; // @[Arbiter.scala 31:68]
  wire  _T_95; // @[Arbiter.scala 31:68]
  wire [29:0] Arbiter_1_covSum;
  assign _GEN_2 = io_in_2_valid ? io_in_2_bits_eccMask : io_in_3_bits_eccMask; // @[Arbiter.scala 126:27]
  assign _GEN_5 = io_in_2_valid ? io_in_2_bits_wdata : io_in_3_bits_wdata; // @[Arbiter.scala 126:27]
  assign _GEN_7 = io_in_2_valid ? io_in_2_bits_addr : io_in_3_bits_addr; // @[Arbiter.scala 126:27]
  assign _GEN_9 = io_in_1_valid ? io_in_1_bits_way_en : 4'hf; // @[Arbiter.scala 126:27]
  assign _GEN_10 = io_in_1_valid ? 8'hff : _GEN_2; // @[Arbiter.scala 126:27]
  assign _GEN_13 = io_in_1_valid ? io_in_1_bits_wdata : _GEN_5; // @[Arbiter.scala 126:27]
  assign _GEN_14 = io_in_1_valid & io_in_1_bits_write; // @[Arbiter.scala 126:27]
  assign _GEN_15 = io_in_1_valid ? io_in_1_bits_addr : _GEN_7; // @[Arbiter.scala 126:27]
  assign _T_94 = io_in_0_valid | io_in_1_valid; // @[Arbiter.scala 31:68]
  assign _T_95 = _T_94 | io_in_2_valid; // @[Arbiter.scala 31:68]
  assign io_in_1_ready = ~io_in_0_valid; // @[Arbiter.scala 134:14]
  assign io_in_2_ready = ~_T_94; // @[Arbiter.scala 134:14]
  assign io_in_3_ready = ~_T_95; // @[Arbiter.scala 134:14]
  assign io_out_valid = _T_95 | io_in_3_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_15; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_write = io_in_0_valid ? io_in_0_bits_write : _GEN_14; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_wdata = io_in_0_valid ? io_in_0_bits_wdata : _GEN_13; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_eccMask = io_in_0_valid ? io_in_0_bits_eccMask : _GEN_10; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_way_en = io_in_0_valid ? io_in_0_bits_way_en : _GEN_9; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign Arbiter_1_covSum = 30'h0;
  assign io_covSum = Arbiter_1_covSum;
  assign metaAssert = 1'h0;
endmodule
module TLB(
  input         clock,
  input         reset,
  output        io_req_ready,
  input         io_req_valid,
  input  [39:0] io_req_bits_vaddr,
  input         io_req_bits_passthrough,
  input  [1:0]  io_req_bits_size,
  input  [4:0]  io_req_bits_cmd,
  output        io_resp_miss,
  output [31:0] io_resp_paddr,
  output        io_resp_pf_ld,
  output        io_resp_pf_st,
  output        io_resp_ae_ld,
  output        io_resp_ae_st,
  output        io_resp_ma_ld,
  output        io_resp_ma_st,
  output        io_resp_cacheable,
  input         io_sfence_valid,
  input         io_sfence_bits_rs1,
  input         io_sfence_bits_rs2,
  input  [38:0] io_sfence_bits_addr,
  input         io_ptw_req_ready,
  output        io_ptw_req_valid,
  output        io_ptw_req_bits_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  input         io_ptw_resp_valid,
  input         io_ptw_resp_bits_ae,
  input  [53:0] io_ptw_resp_bits_pte_ppn,
  input         io_ptw_resp_bits_pte_d,
  input         io_ptw_resp_bits_pte_a,
  input         io_ptw_resp_bits_pte_g,
  input         io_ptw_resp_bits_pte_u,
  input         io_ptw_resp_bits_pte_x,
  input         io_ptw_resp_bits_pte_w,
  input         io_ptw_resp_bits_pte_r,
  input         io_ptw_resp_bits_pte_v,
  input  [1:0]  io_ptw_resp_bits_level,
  input         io_ptw_resp_bits_homogeneous,
  input  [3:0]  io_ptw_ptbr_mode,
  input  [1:0]  io_ptw_status_dprv,
  input         io_ptw_status_mxr,
  input         io_ptw_status_sum,
  input         io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
  input         io_ptw_pmp_0_cfg_w,
  input         io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr,
  input  [31:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
  input         io_ptw_pmp_1_cfg_w,
  input         io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr,
  input  [31:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
  input         io_ptw_pmp_2_cfg_w,
  input         io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr,
  input  [31:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
  input         io_ptw_pmp_3_cfg_w,
  input         io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr,
  input  [31:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
  input         io_ptw_pmp_4_cfg_w,
  input         io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr,
  input  [31:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
  input         io_ptw_pmp_5_cfg_w,
  input         io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr,
  input  [31:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
  input         io_ptw_pmp_6_cfg_w,
  input         io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr,
  input  [31:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
  input         io_ptw_pmp_7_cfg_w,
  input         io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr,
  input  [31:0] io_ptw_pmp_7_mask,
  input  [26:0] io_ptw_vpoffset_bits_value,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [1:0] pmp_io_prv; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_0_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_0_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_0_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_0_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_0_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_0_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_0_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_1_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_1_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_1_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_1_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_1_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_1_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_1_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_2_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_2_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_2_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_2_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_2_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_2_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_2_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_3_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_3_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_3_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_3_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_3_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_3_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_3_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_4_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_4_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_4_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_4_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_4_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_4_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_4_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_5_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_5_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_5_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_5_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_5_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_5_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_5_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_6_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_6_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_6_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_6_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_6_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_6_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_6_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_7_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_7_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_7_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_7_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_7_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_7_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_7_mask; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_addr; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_size; // @[TLB.scala 190:19]
  wire  pmp_io_r; // @[TLB.scala 190:19]
  wire  pmp_io_w; // @[TLB.scala 190:19]
  wire  pmp_io_x; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_covSum; // @[TLB.scala 190:19]
  wire  pmp_metaAssert; // @[TLB.scala 190:19]
  reg [26:0] sectored_entries_0_tag; // @[TLB.scala 163:29]
  reg [31:0] _RAND_0;
  reg [33:0] sectored_entries_0_data_0; // @[TLB.scala 163:29]
  reg [63:0] _RAND_1;
  reg [33:0] sectored_entries_0_data_1; // @[TLB.scala 163:29]
  reg [63:0] _RAND_2;
  reg [33:0] sectored_entries_0_data_2; // @[TLB.scala 163:29]
  reg [63:0] _RAND_3;
  reg [33:0] sectored_entries_0_data_3; // @[TLB.scala 163:29]
  reg [63:0] _RAND_4;
  reg  sectored_entries_0_valid_0; // @[TLB.scala 163:29]
  reg [31:0] _RAND_5;
  reg  sectored_entries_0_valid_1; // @[TLB.scala 163:29]
  reg [31:0] _RAND_6;
  reg  sectored_entries_0_valid_2; // @[TLB.scala 163:29]
  reg [31:0] _RAND_7;
  reg  sectored_entries_0_valid_3; // @[TLB.scala 163:29]
  reg [31:0] _RAND_8;
  reg [26:0] sectored_entries_1_tag; // @[TLB.scala 163:29]
  reg [31:0] _RAND_9;
  reg [33:0] sectored_entries_1_data_0; // @[TLB.scala 163:29]
  reg [63:0] _RAND_10;
  reg [33:0] sectored_entries_1_data_1; // @[TLB.scala 163:29]
  reg [63:0] _RAND_11;
  reg [33:0] sectored_entries_1_data_2; // @[TLB.scala 163:29]
  reg [63:0] _RAND_12;
  reg [33:0] sectored_entries_1_data_3; // @[TLB.scala 163:29]
  reg [63:0] _RAND_13;
  reg  sectored_entries_1_valid_0; // @[TLB.scala 163:29]
  reg [31:0] _RAND_14;
  reg  sectored_entries_1_valid_1; // @[TLB.scala 163:29]
  reg [31:0] _RAND_15;
  reg  sectored_entries_1_valid_2; // @[TLB.scala 163:29]
  reg [31:0] _RAND_16;
  reg  sectored_entries_1_valid_3; // @[TLB.scala 163:29]
  reg [31:0] _RAND_17;
  reg [26:0] sectored_entries_2_tag; // @[TLB.scala 163:29]
  reg [31:0] _RAND_18;
  reg [33:0] sectored_entries_2_data_0; // @[TLB.scala 163:29]
  reg [63:0] _RAND_19;
  reg [33:0] sectored_entries_2_data_1; // @[TLB.scala 163:29]
  reg [63:0] _RAND_20;
  reg [33:0] sectored_entries_2_data_2; // @[TLB.scala 163:29]
  reg [63:0] _RAND_21;
  reg [33:0] sectored_entries_2_data_3; // @[TLB.scala 163:29]
  reg [63:0] _RAND_22;
  reg  sectored_entries_2_valid_0; // @[TLB.scala 163:29]
  reg [31:0] _RAND_23;
  reg  sectored_entries_2_valid_1; // @[TLB.scala 163:29]
  reg [31:0] _RAND_24;
  reg  sectored_entries_2_valid_2; // @[TLB.scala 163:29]
  reg [31:0] _RAND_25;
  reg  sectored_entries_2_valid_3; // @[TLB.scala 163:29]
  reg [31:0] _RAND_26;
  reg [26:0] sectored_entries_3_tag; // @[TLB.scala 163:29]
  reg [31:0] _RAND_27;
  reg [33:0] sectored_entries_3_data_0; // @[TLB.scala 163:29]
  reg [63:0] _RAND_28;
  reg [33:0] sectored_entries_3_data_1; // @[TLB.scala 163:29]
  reg [63:0] _RAND_29;
  reg [33:0] sectored_entries_3_data_2; // @[TLB.scala 163:29]
  reg [63:0] _RAND_30;
  reg [33:0] sectored_entries_3_data_3; // @[TLB.scala 163:29]
  reg [63:0] _RAND_31;
  reg  sectored_entries_3_valid_0; // @[TLB.scala 163:29]
  reg [31:0] _RAND_32;
  reg  sectored_entries_3_valid_1; // @[TLB.scala 163:29]
  reg [31:0] _RAND_33;
  reg  sectored_entries_3_valid_2; // @[TLB.scala 163:29]
  reg [31:0] _RAND_34;
  reg  sectored_entries_3_valid_3; // @[TLB.scala 163:29]
  reg [31:0] _RAND_35;
  reg [26:0] sectored_entries_4_tag; // @[TLB.scala 163:29]
  reg [31:0] _RAND_36;
  reg [33:0] sectored_entries_4_data_0; // @[TLB.scala 163:29]
  reg [63:0] _RAND_37;
  reg [33:0] sectored_entries_4_data_1; // @[TLB.scala 163:29]
  reg [63:0] _RAND_38;
  reg [33:0] sectored_entries_4_data_2; // @[TLB.scala 163:29]
  reg [63:0] _RAND_39;
  reg [33:0] sectored_entries_4_data_3; // @[TLB.scala 163:29]
  reg [63:0] _RAND_40;
  reg  sectored_entries_4_valid_0; // @[TLB.scala 163:29]
  reg [31:0] _RAND_41;
  reg  sectored_entries_4_valid_1; // @[TLB.scala 163:29]
  reg [31:0] _RAND_42;
  reg  sectored_entries_4_valid_2; // @[TLB.scala 163:29]
  reg [31:0] _RAND_43;
  reg  sectored_entries_4_valid_3; // @[TLB.scala 163:29]
  reg [31:0] _RAND_44;
  reg [26:0] sectored_entries_5_tag; // @[TLB.scala 163:29]
  reg [31:0] _RAND_45;
  reg [33:0] sectored_entries_5_data_0; // @[TLB.scala 163:29]
  reg [63:0] _RAND_46;
  reg [33:0] sectored_entries_5_data_1; // @[TLB.scala 163:29]
  reg [63:0] _RAND_47;
  reg [33:0] sectored_entries_5_data_2; // @[TLB.scala 163:29]
  reg [63:0] _RAND_48;
  reg [33:0] sectored_entries_5_data_3; // @[TLB.scala 163:29]
  reg [63:0] _RAND_49;
  reg  sectored_entries_5_valid_0; // @[TLB.scala 163:29]
  reg [31:0] _RAND_50;
  reg  sectored_entries_5_valid_1; // @[TLB.scala 163:29]
  reg [31:0] _RAND_51;
  reg  sectored_entries_5_valid_2; // @[TLB.scala 163:29]
  reg [31:0] _RAND_52;
  reg  sectored_entries_5_valid_3; // @[TLB.scala 163:29]
  reg [31:0] _RAND_53;
  reg [26:0] sectored_entries_6_tag; // @[TLB.scala 163:29]
  reg [31:0] _RAND_54;
  reg [33:0] sectored_entries_6_data_0; // @[TLB.scala 163:29]
  reg [63:0] _RAND_55;
  reg [33:0] sectored_entries_6_data_1; // @[TLB.scala 163:29]
  reg [63:0] _RAND_56;
  reg [33:0] sectored_entries_6_data_2; // @[TLB.scala 163:29]
  reg [63:0] _RAND_57;
  reg [33:0] sectored_entries_6_data_3; // @[TLB.scala 163:29]
  reg [63:0] _RAND_58;
  reg  sectored_entries_6_valid_0; // @[TLB.scala 163:29]
  reg [31:0] _RAND_59;
  reg  sectored_entries_6_valid_1; // @[TLB.scala 163:29]
  reg [31:0] _RAND_60;
  reg  sectored_entries_6_valid_2; // @[TLB.scala 163:29]
  reg [31:0] _RAND_61;
  reg  sectored_entries_6_valid_3; // @[TLB.scala 163:29]
  reg [31:0] _RAND_62;
  reg [26:0] sectored_entries_7_tag; // @[TLB.scala 163:29]
  reg [31:0] _RAND_63;
  reg [33:0] sectored_entries_7_data_0; // @[TLB.scala 163:29]
  reg [63:0] _RAND_64;
  reg [33:0] sectored_entries_7_data_1; // @[TLB.scala 163:29]
  reg [63:0] _RAND_65;
  reg [33:0] sectored_entries_7_data_2; // @[TLB.scala 163:29]
  reg [63:0] _RAND_66;
  reg [33:0] sectored_entries_7_data_3; // @[TLB.scala 163:29]
  reg [63:0] _RAND_67;
  reg  sectored_entries_7_valid_0; // @[TLB.scala 163:29]
  reg [31:0] _RAND_68;
  reg  sectored_entries_7_valid_1; // @[TLB.scala 163:29]
  reg [31:0] _RAND_69;
  reg  sectored_entries_7_valid_2; // @[TLB.scala 163:29]
  reg [31:0] _RAND_70;
  reg  sectored_entries_7_valid_3; // @[TLB.scala 163:29]
  reg [31:0] _RAND_71;
  reg [1:0] superpage_entries_0_level; // @[TLB.scala 164:30]
  reg [31:0] _RAND_72;
  reg [26:0] superpage_entries_0_tag; // @[TLB.scala 164:30]
  reg [31:0] _RAND_73;
  reg [33:0] superpage_entries_0_data_0; // @[TLB.scala 164:30]
  reg [63:0] _RAND_74;
  reg  superpage_entries_0_valid_0; // @[TLB.scala 164:30]
  reg [31:0] _RAND_75;
  reg [1:0] superpage_entries_1_level; // @[TLB.scala 164:30]
  reg [31:0] _RAND_76;
  reg [26:0] superpage_entries_1_tag; // @[TLB.scala 164:30]
  reg [31:0] _RAND_77;
  reg [33:0] superpage_entries_1_data_0; // @[TLB.scala 164:30]
  reg [63:0] _RAND_78;
  reg  superpage_entries_1_valid_0; // @[TLB.scala 164:30]
  reg [31:0] _RAND_79;
  reg [1:0] superpage_entries_2_level; // @[TLB.scala 164:30]
  reg [31:0] _RAND_80;
  reg [26:0] superpage_entries_2_tag; // @[TLB.scala 164:30]
  reg [31:0] _RAND_81;
  reg [33:0] superpage_entries_2_data_0; // @[TLB.scala 164:30]
  reg [63:0] _RAND_82;
  reg  superpage_entries_2_valid_0; // @[TLB.scala 164:30]
  reg [31:0] _RAND_83;
  reg [1:0] superpage_entries_3_level; // @[TLB.scala 164:30]
  reg [31:0] _RAND_84;
  reg [26:0] superpage_entries_3_tag; // @[TLB.scala 164:30]
  reg [31:0] _RAND_85;
  reg [33:0] superpage_entries_3_data_0; // @[TLB.scala 164:30]
  reg [63:0] _RAND_86;
  reg  superpage_entries_3_valid_0; // @[TLB.scala 164:30]
  reg [31:0] _RAND_87;
  reg [1:0] special_entry_level; // @[TLB.scala 165:56]
  reg [31:0] _RAND_88;
  reg [26:0] special_entry_tag; // @[TLB.scala 165:56]
  reg [31:0] _RAND_89;
  reg [33:0] special_entry_data_0; // @[TLB.scala 165:56]
  reg [63:0] _RAND_90;
  reg  special_entry_valid_0; // @[TLB.scala 165:56]
  reg [31:0] _RAND_91;
  reg [1:0] state; // @[TLB.scala 170:18]
  reg [31:0] _RAND_92;
  reg [26:0] r_refill_tag; // @[TLB.scala 171:25]
  reg [31:0] _RAND_93;
  reg [1:0] r_superpage_repl_addr; // @[TLB.scala 172:34]
  reg [31:0] _RAND_94;
  reg [2:0] r_sectored_repl_addr; // @[TLB.scala 173:33]
  reg [31:0] _RAND_95;
  reg [2:0] r_sectored_hit_addr; // @[TLB.scala 174:32]
  reg [31:0] _RAND_96;
  reg  r_sectored_hit; // @[TLB.scala 175:27]
  reg [31:0] _RAND_97;
  wire  priv_s; // @[TLB.scala 178:20]
  wire  priv_uses_vm; // @[TLB.scala 179:27]
  wire  _T_322; // @[TLB.scala 180:83]
  wire  vm_enabled; // @[TLB.scala 180:99]
  wire [26:0] vpn; // @[TLB.scala 183:30]
  wire [19:0] refill_ppn; // @[TLB.scala 184:44]
  wire  _T_324; // @[package.scala 14:47]
  wire  _T_325; // @[package.scala 14:47]
  wire  invalidate_refill; // @[package.scala 14:62]
  wire  _T_348; // @[TLB.scala 123:30]
  wire [26:0] _T_350; // @[TLB.scala 124:30]
  wire [26:0] _GEN_954; // @[TLB.scala 124:49]
  wire [26:0] _T_351; // @[TLB.scala 124:49]
  wire  _T_354; // @[TLB.scala 123:30]
  wire [26:0] _T_356; // @[TLB.scala 124:30]
  wire [26:0] _T_357; // @[TLB.scala 124:49]
  wire [19:0] _T_359; // @[Cat.scala 30:58]
  wire [27:0] _T_361; // @[TLB.scala 188:20]
  wire [27:0] mpu_ppn; // @[TLB.scala 187:20]
  wire [39:0] mpu_physaddr; // @[Cat.scala 30:58]
  wire  _T_363; // @[TLB.scala 194:49]
  wire [39:0] _T_366; // @[Parameters.scala 121:31]
  wire [40:0] _T_367; // @[Parameters.scala 121:49]
  wire [40:0] _T_369; // @[Parameters.scala 121:52]
  wire  _T_370; // @[Parameters.scala 121:67]
  wire [39:0] _T_371; // @[Parameters.scala 121:31]
  wire [40:0] _T_372; // @[Parameters.scala 121:49]
  wire [40:0] _T_374; // @[Parameters.scala 121:52]
  wire  _T_375; // @[Parameters.scala 121:67]
  wire [39:0] _T_376; // @[Parameters.scala 121:31]
  wire [40:0] _T_377; // @[Parameters.scala 121:49]
  wire [40:0] _T_379; // @[Parameters.scala 121:52]
  wire  _T_380; // @[Parameters.scala 121:67]
  wire [40:0] _T_382; // @[Parameters.scala 121:49]
  wire [40:0] _T_384; // @[Parameters.scala 121:52]
  wire  _T_385; // @[Parameters.scala 121:67]
  wire [39:0] _T_386; // @[Parameters.scala 121:31]
  wire [40:0] _T_387; // @[Parameters.scala 121:49]
  wire [40:0] _T_389; // @[Parameters.scala 121:52]
  wire  _T_390; // @[Parameters.scala 121:67]
  wire [39:0] _T_391; // @[Parameters.scala 121:31]
  wire [40:0] _T_392; // @[Parameters.scala 121:49]
  wire [40:0] _T_394; // @[Parameters.scala 121:52]
  wire  _T_395; // @[Parameters.scala 121:67]
  wire [39:0] _T_396; // @[Parameters.scala 121:31]
  wire [40:0] _T_397; // @[Parameters.scala 121:49]
  wire [40:0] _T_399; // @[Parameters.scala 121:52]
  wire  _T_400; // @[Parameters.scala 121:67]
  wire  _T_414; // @[TLB.scala 195:67]
  wire  _T_415; // @[TLB.scala 195:67]
  wire  _T_416; // @[TLB.scala 195:67]
  wire  _T_417; // @[TLB.scala 195:67]
  wire  _T_418; // @[TLB.scala 195:67]
  wire  legal_address; // @[TLB.scala 195:67]
  wire [40:0] _T_427; // @[Parameters.scala 121:52]
  wire  _T_428; // @[Parameters.scala 121:67]
  wire  cacheable; // @[TLB.scala 197:19]
  wire [39:0] _T_485; // @[Parameters.scala 121:31]
  wire [40:0] _T_486; // @[Parameters.scala 121:49]
  wire [40:0] _T_488; // @[Parameters.scala 121:52]
  wire  _T_489; // @[Parameters.scala 121:67]
  wire [40:0] _T_507; // @[Parameters.scala 121:52]
  wire  _T_508; // @[Parameters.scala 121:67]
  wire  _T_515; // @[TLBPermissions.scala 81:66]
  wire  prot_r; // @[TLB.scala 200:41]
  wire [40:0] _T_552; // @[Parameters.scala 121:52]
  wire  _T_553; // @[Parameters.scala 121:67]
  wire [39:0] _T_554; // @[Parameters.scala 121:31]
  wire [40:0] _T_555; // @[Parameters.scala 121:49]
  wire [40:0] _T_557; // @[Parameters.scala 121:52]
  wire  _T_558; // @[Parameters.scala 121:67]
  wire  _T_560; // @[Parameters.scala 148:89]
  wire  _T_561; // @[Parameters.scala 148:89]
  wire  _T_568; // @[TLB.scala 197:19]
  wire  prot_w; // @[TLB.scala 201:45]
  wire  _T_603; // @[TLB.scala 197:19]
  wire  prot_al; // @[TLB.scala 202:46]
  wire [40:0] _T_655; // @[Parameters.scala 121:52]
  wire  _T_656; // @[Parameters.scala 121:67]
  wire  _T_667; // @[Parameters.scala 148:89]
  wire  _T_668; // @[Parameters.scala 148:89]
  wire  _T_675; // @[TLB.scala 197:19]
  wire  prot_x; // @[TLB.scala 204:40]
  wire [40:0] _T_701; // @[Parameters.scala 121:52]
  wire  _T_702; // @[Parameters.scala 121:67]
  wire [40:0] _T_706; // @[Parameters.scala 121:52]
  wire  _T_707; // @[Parameters.scala 121:67]
  wire  _T_713; // @[Parameters.scala 148:89]
  wire  _T_714; // @[Parameters.scala 148:89]
  wire  _T_715; // @[Parameters.scala 148:89]
  wire  prot_eff; // @[TLB.scala 197:19]
  wire  _T_722; // @[package.scala 63:59]
  wire  _T_723; // @[package.scala 63:59]
  wire  _T_724; // @[package.scala 63:59]
  wire [26:0] _T_725; // @[TLB.scala 103:43]
  wire  _T_727; // @[TLB.scala 103:68]
  wire  sector_hits_0; // @[TLB.scala 102:42]
  wire  _T_728; // @[package.scala 63:59]
  wire  _T_729; // @[package.scala 63:59]
  wire  _T_730; // @[package.scala 63:59]
  wire [26:0] _T_731; // @[TLB.scala 103:43]
  wire  _T_733; // @[TLB.scala 103:68]
  wire  sector_hits_1; // @[TLB.scala 102:42]
  wire  _T_734; // @[package.scala 63:59]
  wire  _T_735; // @[package.scala 63:59]
  wire  _T_736; // @[package.scala 63:59]
  wire [26:0] _T_737; // @[TLB.scala 103:43]
  wire  _T_739; // @[TLB.scala 103:68]
  wire  sector_hits_2; // @[TLB.scala 102:42]
  wire  _T_740; // @[package.scala 63:59]
  wire  _T_741; // @[package.scala 63:59]
  wire  _T_742; // @[package.scala 63:59]
  wire [26:0] _T_743; // @[TLB.scala 103:43]
  wire  _T_745; // @[TLB.scala 103:68]
  wire  sector_hits_3; // @[TLB.scala 102:42]
  wire  _T_746; // @[package.scala 63:59]
  wire  _T_747; // @[package.scala 63:59]
  wire  _T_748; // @[package.scala 63:59]
  wire [26:0] _T_749; // @[TLB.scala 103:43]
  wire  _T_751; // @[TLB.scala 103:68]
  wire  sector_hits_4; // @[TLB.scala 102:42]
  wire  _T_752; // @[package.scala 63:59]
  wire  _T_753; // @[package.scala 63:59]
  wire  _T_754; // @[package.scala 63:59]
  wire [26:0] _T_755; // @[TLB.scala 103:43]
  wire  _T_757; // @[TLB.scala 103:68]
  wire  sector_hits_5; // @[TLB.scala 102:42]
  wire  _T_758; // @[package.scala 63:59]
  wire  _T_759; // @[package.scala 63:59]
  wire  _T_760; // @[package.scala 63:59]
  wire [26:0] _T_761; // @[TLB.scala 103:43]
  wire  _T_763; // @[TLB.scala 103:68]
  wire  sector_hits_6; // @[TLB.scala 102:42]
  wire  _T_764; // @[package.scala 63:59]
  wire  _T_765; // @[package.scala 63:59]
  wire  _T_766; // @[package.scala 63:59]
  wire [26:0] _T_767; // @[TLB.scala 103:43]
  wire  _T_769; // @[TLB.scala 103:68]
  wire  sector_hits_7; // @[TLB.scala 102:42]
  wire  _T_774; // @[TLB.scala 110:79]
  wire  _T_776; // @[TLB.scala 110:31]
  wire  _T_777; // @[TLB.scala 109:30]
  wire  _T_781; // @[TLB.scala 110:79]
  wire  _T_782; // @[TLB.scala 110:42]
  wire  superpage_hits_0; // @[TLB.scala 110:31]
  wire  _T_794; // @[TLB.scala 110:79]
  wire  _T_796; // @[TLB.scala 110:31]
  wire  _T_797; // @[TLB.scala 109:30]
  wire  _T_801; // @[TLB.scala 110:79]
  wire  _T_802; // @[TLB.scala 110:42]
  wire  superpage_hits_1; // @[TLB.scala 110:31]
  wire  _T_814; // @[TLB.scala 110:79]
  wire  _T_816; // @[TLB.scala 110:31]
  wire  _T_817; // @[TLB.scala 109:30]
  wire  _T_821; // @[TLB.scala 110:79]
  wire  _T_822; // @[TLB.scala 110:42]
  wire  superpage_hits_2; // @[TLB.scala 110:31]
  wire  _T_834; // @[TLB.scala 110:79]
  wire  _T_836; // @[TLB.scala 110:31]
  wire  _T_837; // @[TLB.scala 109:30]
  wire  _T_841; // @[TLB.scala 110:79]
  wire  _T_842; // @[TLB.scala 110:42]
  wire  superpage_hits_3; // @[TLB.scala 110:31]
  wire  _GEN_1; // @[TLB.scala 115:20]
  wire  _GEN_2; // @[TLB.scala 115:20]
  wire  _GEN_3; // @[TLB.scala 115:20]
  wire  _T_854; // @[TLB.scala 115:20]
  wire  hitsVec_0; // @[TLB.scala 209:44]
  wire  _GEN_5; // @[TLB.scala 115:20]
  wire  _GEN_6; // @[TLB.scala 115:20]
  wire  _GEN_7; // @[TLB.scala 115:20]
  wire  _T_859; // @[TLB.scala 115:20]
  wire  hitsVec_1; // @[TLB.scala 209:44]
  wire  _GEN_9; // @[TLB.scala 115:20]
  wire  _GEN_10; // @[TLB.scala 115:20]
  wire  _GEN_11; // @[TLB.scala 115:20]
  wire  _T_864; // @[TLB.scala 115:20]
  wire  hitsVec_2; // @[TLB.scala 209:44]
  wire  _GEN_13; // @[TLB.scala 115:20]
  wire  _GEN_14; // @[TLB.scala 115:20]
  wire  _GEN_15; // @[TLB.scala 115:20]
  wire  _T_869; // @[TLB.scala 115:20]
  wire  hitsVec_3; // @[TLB.scala 209:44]
  wire  _GEN_17; // @[TLB.scala 115:20]
  wire  _GEN_18; // @[TLB.scala 115:20]
  wire  _GEN_19; // @[TLB.scala 115:20]
  wire  _T_874; // @[TLB.scala 115:20]
  wire  hitsVec_4; // @[TLB.scala 209:44]
  wire  _GEN_21; // @[TLB.scala 115:20]
  wire  _GEN_22; // @[TLB.scala 115:20]
  wire  _GEN_23; // @[TLB.scala 115:20]
  wire  _T_879; // @[TLB.scala 115:20]
  wire  hitsVec_5; // @[TLB.scala 209:44]
  wire  _GEN_25; // @[TLB.scala 115:20]
  wire  _GEN_26; // @[TLB.scala 115:20]
  wire  _GEN_27; // @[TLB.scala 115:20]
  wire  _T_884; // @[TLB.scala 115:20]
  wire  hitsVec_6; // @[TLB.scala 209:44]
  wire  _GEN_29; // @[TLB.scala 115:20]
  wire  _GEN_30; // @[TLB.scala 115:20]
  wire  _GEN_31; // @[TLB.scala 115:20]
  wire  _T_889; // @[TLB.scala 115:20]
  wire  hitsVec_7; // @[TLB.scala 209:44]
  wire  hitsVec_8; // @[TLB.scala 209:44]
  wire  hitsVec_9; // @[TLB.scala 209:44]
  wire  hitsVec_10; // @[TLB.scala 209:44]
  wire  hitsVec_11; // @[TLB.scala 209:44]
  wire  _T_978; // @[TLB.scala 110:79]
  wire  _T_980; // @[TLB.scala 110:31]
  wire  _T_985; // @[TLB.scala 110:79]
  wire  _T_986; // @[TLB.scala 110:42]
  wire  _T_987; // @[TLB.scala 110:31]
  wire  _T_992; // @[TLB.scala 110:79]
  wire  _T_993; // @[TLB.scala 110:42]
  wire  _T_994; // @[TLB.scala 110:31]
  wire  hitsVec_12; // @[TLB.scala 209:44]
  wire [5:0] _T_999; // @[Cat.scala 30:58]
  wire [12:0] real_hits; // @[Cat.scala 30:58]
  wire [13:0] hits; // @[Cat.scala 30:58]
  wire [33:0] _GEN_33;
  wire [33:0] _GEN_34;
  wire [33:0] _GEN_35;
  wire [33:0] _GEN_37;
  wire [33:0] _GEN_38;
  wire [33:0] _GEN_39;
  wire [33:0] _GEN_41;
  wire [33:0] _GEN_42;
  wire [33:0] _GEN_43;
  wire [33:0] _GEN_45;
  wire [33:0] _GEN_46;
  wire [33:0] _GEN_47;
  wire [33:0] _GEN_49;
  wire [33:0] _GEN_50;
  wire [33:0] _GEN_51;
  wire [33:0] _GEN_53;
  wire [33:0] _GEN_54;
  wire [33:0] _GEN_55;
  wire [33:0] _GEN_57;
  wire [33:0] _GEN_58;
  wire [33:0] _GEN_59;
  wire [33:0] _GEN_61;
  wire [33:0] _GEN_62;
  wire [33:0] _GEN_63;
  wire [26:0] _T_1199; // @[TLB.scala 124:30]
  wire [26:0] _GEN_956; // @[TLB.scala 124:49]
  wire [26:0] _T_1200; // @[TLB.scala 124:49]
  wire [26:0] _T_1206; // @[TLB.scala 124:49]
  wire [19:0] _T_1208; // @[Cat.scala 30:58]
  wire [26:0] _T_1232; // @[TLB.scala 124:30]
  wire [26:0] _GEN_958; // @[TLB.scala 124:49]
  wire [26:0] _T_1233; // @[TLB.scala 124:49]
  wire [26:0] _T_1239; // @[TLB.scala 124:49]
  wire [19:0] _T_1241; // @[Cat.scala 30:58]
  wire [26:0] _T_1265; // @[TLB.scala 124:30]
  wire [26:0] _GEN_960; // @[TLB.scala 124:49]
  wire [26:0] _T_1266; // @[TLB.scala 124:49]
  wire [26:0] _T_1272; // @[TLB.scala 124:49]
  wire [19:0] _T_1274; // @[Cat.scala 30:58]
  wire [26:0] _T_1298; // @[TLB.scala 124:30]
  wire [26:0] _GEN_962; // @[TLB.scala 124:49]
  wire [26:0] _T_1299; // @[TLB.scala 124:49]
  wire [26:0] _T_1305; // @[TLB.scala 124:49]
  wire [19:0] _T_1307; // @[Cat.scala 30:58]
  wire [19:0] _T_1343; // @[Mux.scala 19:72]
  wire [19:0] _T_1344; // @[Mux.scala 19:72]
  wire [19:0] _T_1345; // @[Mux.scala 19:72]
  wire [19:0] _T_1346; // @[Mux.scala 19:72]
  wire [19:0] _T_1347; // @[Mux.scala 19:72]
  wire [19:0] _T_1348; // @[Mux.scala 19:72]
  wire [19:0] _T_1349; // @[Mux.scala 19:72]
  wire [19:0] _T_1350; // @[Mux.scala 19:72]
  wire [19:0] _T_1351; // @[Mux.scala 19:72]
  wire [19:0] _T_1352; // @[Mux.scala 19:72]
  wire [19:0] _T_1353; // @[Mux.scala 19:72]
  wire [19:0] _T_1354; // @[Mux.scala 19:72]
  wire [19:0] _T_1355; // @[Mux.scala 19:72]
  wire [19:0] _T_1356; // @[Mux.scala 19:72]
  wire [19:0] _T_1357; // @[Mux.scala 19:72]
  wire [19:0] _T_1358; // @[Mux.scala 19:72]
  wire [19:0] _T_1359; // @[Mux.scala 19:72]
  wire [19:0] _T_1360; // @[Mux.scala 19:72]
  wire [19:0] _T_1361; // @[Mux.scala 19:72]
  wire [19:0] _T_1362; // @[Mux.scala 19:72]
  wire [19:0] _T_1363; // @[Mux.scala 19:72]
  wire [19:0] _T_1364; // @[Mux.scala 19:72]
  wire [19:0] _T_1365; // @[Mux.scala 19:72]
  wire [19:0] _T_1366; // @[Mux.scala 19:72]
  wire [19:0] _T_1367; // @[Mux.scala 19:72]
  wire [19:0] _T_1368; // @[Mux.scala 19:72]
  wire [19:0] ppn; // @[Mux.scala 19:72]
  reg [26:0] vpoffset_cfg_value; // @[TLB.scala 215:29]
  reg [31:0] _RAND_98;
  reg [26:0] requestedVPN; // @[TLB.scala 216:25]
  reg [31:0] _RAND_99;
  wire  _T_1385; // @[TLB.scala 224:17]
  wire [53:0] _GEN_966; // @[TLB.scala 227:31]
  wire [53:0] _T_1387; // @[TLB.scala 227:31]
  wire  _T_1391; // @[PTW.scala 77:44]
  wire  _T_1392; // @[PTW.scala 77:38]
  wire  _T_1393; // @[PTW.scala 77:32]
  wire  _T_1394; // @[PTW.scala 77:52]
  wire  _T_1395; // @[PTW.scala 81:35]
  wire  _T_1401; // @[PTW.scala 82:35]
  wire  _T_1402; // @[PTW.scala 82:40]
  wire  _T_1403; // @[TLB.scala 231:55]
  wire  _T_1404; // @[TLB.scala 231:32]
  wire  _T_1405; // @[TLB.scala 231:90]
  wire  _T_1406; // @[TLB.scala 231:64]
  wire  _T_1412; // @[PTW.scala 83:35]
  wire [53:0] _GEN_967; // @[TLB.scala 231:133]
  wire  _T_1413; // @[TLB.scala 231:133]
  wire  _T_1420; // @[TLB.scala 231:120]
  wire  _T_1421; // @[TLB.scala 231:25]
  wire [6:0] _T_1430; // @[TLB.scala 138:26]
  wire [33:0] _T_1438; // @[TLB.scala 138:26]
  wire  _T_1439; // @[TLB.scala 253:40]
  wire  _T_1440; // @[TLB.scala 254:82]
  wire  _GEN_67; // @[TLB.scala 254:89]
  wire  _T_1456; // @[TLB.scala 254:82]
  wire  _GEN_71; // @[TLB.scala 254:89]
  wire  _T_1472; // @[TLB.scala 254:82]
  wire  _GEN_75; // @[TLB.scala 254:89]
  wire  _T_1488; // @[TLB.scala 254:82]
  wire  _GEN_79; // @[TLB.scala 254:89]
  wire [2:0] _T_1504; // @[TLB.scala 258:22]
  wire  _T_1505; // @[TLB.scala 259:65]
  wire  _GEN_81; // @[TLB.scala 260:32]
  wire  _GEN_82; // @[TLB.scala 260:32]
  wire  _GEN_83; // @[TLB.scala 260:32]
  wire  _GEN_84; // @[TLB.scala 260:32]
  wire  _GEN_968; // @[TLB.scala 137:18]
  wire  _GEN_85; // @[TLB.scala 137:18]
  wire  _GEN_969; // @[TLB.scala 137:18]
  wire  _GEN_86; // @[TLB.scala 137:18]
  wire  _GEN_970; // @[TLB.scala 137:18]
  wire  _GEN_87; // @[TLB.scala 137:18]
  wire  _GEN_971; // @[TLB.scala 137:18]
  wire  _GEN_88; // @[TLB.scala 137:18]
  wire  _GEN_93; // @[TLB.scala 259:72]
  wire  _GEN_94; // @[TLB.scala 259:72]
  wire  _GEN_95; // @[TLB.scala 259:72]
  wire  _GEN_96; // @[TLB.scala 259:72]
  wire  _T_1522; // @[TLB.scala 259:65]
  wire  _GEN_103; // @[TLB.scala 260:32]
  wire  _GEN_104; // @[TLB.scala 260:32]
  wire  _GEN_105; // @[TLB.scala 260:32]
  wire  _GEN_106; // @[TLB.scala 260:32]
  wire  _GEN_107; // @[TLB.scala 137:18]
  wire  _GEN_108; // @[TLB.scala 137:18]
  wire  _GEN_109; // @[TLB.scala 137:18]
  wire  _GEN_110; // @[TLB.scala 137:18]
  wire  _GEN_115; // @[TLB.scala 259:72]
  wire  _GEN_116; // @[TLB.scala 259:72]
  wire  _GEN_117; // @[TLB.scala 259:72]
  wire  _GEN_118; // @[TLB.scala 259:72]
  wire  _T_1539; // @[TLB.scala 259:65]
  wire  _GEN_125; // @[TLB.scala 260:32]
  wire  _GEN_126; // @[TLB.scala 260:32]
  wire  _GEN_127; // @[TLB.scala 260:32]
  wire  _GEN_128; // @[TLB.scala 260:32]
  wire  _GEN_129; // @[TLB.scala 137:18]
  wire  _GEN_130; // @[TLB.scala 137:18]
  wire  _GEN_131; // @[TLB.scala 137:18]
  wire  _GEN_132; // @[TLB.scala 137:18]
  wire  _GEN_137; // @[TLB.scala 259:72]
  wire  _GEN_138; // @[TLB.scala 259:72]
  wire  _GEN_139; // @[TLB.scala 259:72]
  wire  _GEN_140; // @[TLB.scala 259:72]
  wire  _T_1556; // @[TLB.scala 259:65]
  wire  _GEN_147; // @[TLB.scala 260:32]
  wire  _GEN_148; // @[TLB.scala 260:32]
  wire  _GEN_149; // @[TLB.scala 260:32]
  wire  _GEN_150; // @[TLB.scala 260:32]
  wire  _GEN_151; // @[TLB.scala 137:18]
  wire  _GEN_152; // @[TLB.scala 137:18]
  wire  _GEN_153; // @[TLB.scala 137:18]
  wire  _GEN_154; // @[TLB.scala 137:18]
  wire  _GEN_159; // @[TLB.scala 259:72]
  wire  _GEN_160; // @[TLB.scala 259:72]
  wire  _GEN_161; // @[TLB.scala 259:72]
  wire  _GEN_162; // @[TLB.scala 259:72]
  wire  _T_1573; // @[TLB.scala 259:65]
  wire  _GEN_169; // @[TLB.scala 260:32]
  wire  _GEN_170; // @[TLB.scala 260:32]
  wire  _GEN_171; // @[TLB.scala 260:32]
  wire  _GEN_172; // @[TLB.scala 260:32]
  wire  _GEN_173; // @[TLB.scala 137:18]
  wire  _GEN_174; // @[TLB.scala 137:18]
  wire  _GEN_175; // @[TLB.scala 137:18]
  wire  _GEN_176; // @[TLB.scala 137:18]
  wire  _GEN_181; // @[TLB.scala 259:72]
  wire  _GEN_182; // @[TLB.scala 259:72]
  wire  _GEN_183; // @[TLB.scala 259:72]
  wire  _GEN_184; // @[TLB.scala 259:72]
  wire  _T_1590; // @[TLB.scala 259:65]
  wire  _GEN_191; // @[TLB.scala 260:32]
  wire  _GEN_192; // @[TLB.scala 260:32]
  wire  _GEN_193; // @[TLB.scala 260:32]
  wire  _GEN_194; // @[TLB.scala 260:32]
  wire  _GEN_195; // @[TLB.scala 137:18]
  wire  _GEN_196; // @[TLB.scala 137:18]
  wire  _GEN_197; // @[TLB.scala 137:18]
  wire  _GEN_198; // @[TLB.scala 137:18]
  wire  _GEN_203; // @[TLB.scala 259:72]
  wire  _GEN_204; // @[TLB.scala 259:72]
  wire  _GEN_205; // @[TLB.scala 259:72]
  wire  _GEN_206; // @[TLB.scala 259:72]
  wire  _T_1607; // @[TLB.scala 259:65]
  wire  _GEN_213; // @[TLB.scala 260:32]
  wire  _GEN_214; // @[TLB.scala 260:32]
  wire  _GEN_215; // @[TLB.scala 260:32]
  wire  _GEN_216; // @[TLB.scala 260:32]
  wire  _GEN_217; // @[TLB.scala 137:18]
  wire  _GEN_218; // @[TLB.scala 137:18]
  wire  _GEN_219; // @[TLB.scala 137:18]
  wire  _GEN_220; // @[TLB.scala 137:18]
  wire  _GEN_225; // @[TLB.scala 259:72]
  wire  _GEN_226; // @[TLB.scala 259:72]
  wire  _GEN_227; // @[TLB.scala 259:72]
  wire  _GEN_228; // @[TLB.scala 259:72]
  wire  _T_1624; // @[TLB.scala 259:65]
  wire  _GEN_235; // @[TLB.scala 260:32]
  wire  _GEN_236; // @[TLB.scala 260:32]
  wire  _GEN_237; // @[TLB.scala 260:32]
  wire  _GEN_238; // @[TLB.scala 260:32]
  wire  _GEN_239; // @[TLB.scala 137:18]
  wire  _GEN_240; // @[TLB.scala 137:18]
  wire  _GEN_241; // @[TLB.scala 137:18]
  wire  _GEN_242; // @[TLB.scala 137:18]
  wire  _GEN_247; // @[TLB.scala 259:72]
  wire  _GEN_248; // @[TLB.scala 259:72]
  wire  _GEN_249; // @[TLB.scala 259:72]
  wire  _GEN_250; // @[TLB.scala 259:72]
  wire  _GEN_259; // @[TLB.scala 253:54]
  wire  _GEN_263; // @[TLB.scala 253:54]
  wire  _GEN_267; // @[TLB.scala 253:54]
  wire  _GEN_271; // @[TLB.scala 253:54]
  wire  _GEN_273; // @[TLB.scala 253:54]
  wire  _GEN_274; // @[TLB.scala 253:54]
  wire  _GEN_275; // @[TLB.scala 253:54]
  wire  _GEN_276; // @[TLB.scala 253:54]
  wire  _GEN_283; // @[TLB.scala 253:54]
  wire  _GEN_284; // @[TLB.scala 253:54]
  wire  _GEN_285; // @[TLB.scala 253:54]
  wire  _GEN_286; // @[TLB.scala 253:54]
  wire  _GEN_293; // @[TLB.scala 253:54]
  wire  _GEN_294; // @[TLB.scala 253:54]
  wire  _GEN_295; // @[TLB.scala 253:54]
  wire  _GEN_296; // @[TLB.scala 253:54]
  wire  _GEN_303; // @[TLB.scala 253:54]
  wire  _GEN_304; // @[TLB.scala 253:54]
  wire  _GEN_305; // @[TLB.scala 253:54]
  wire  _GEN_306; // @[TLB.scala 253:54]
  wire  _GEN_313; // @[TLB.scala 253:54]
  wire  _GEN_314; // @[TLB.scala 253:54]
  wire  _GEN_315; // @[TLB.scala 253:54]
  wire  _GEN_316; // @[TLB.scala 253:54]
  wire  _GEN_323; // @[TLB.scala 253:54]
  wire  _GEN_324; // @[TLB.scala 253:54]
  wire  _GEN_325; // @[TLB.scala 253:54]
  wire  _GEN_326; // @[TLB.scala 253:54]
  wire  _GEN_333; // @[TLB.scala 253:54]
  wire  _GEN_334; // @[TLB.scala 253:54]
  wire  _GEN_335; // @[TLB.scala 253:54]
  wire  _GEN_336; // @[TLB.scala 253:54]
  wire  _GEN_343; // @[TLB.scala 253:54]
  wire  _GEN_344; // @[TLB.scala 253:54]
  wire  _GEN_345; // @[TLB.scala 253:54]
  wire  _GEN_346; // @[TLB.scala 253:54]
  wire  _GEN_355; // @[TLB.scala 251:68]
  wire  _GEN_359; // @[TLB.scala 251:68]
  wire  _GEN_363; // @[TLB.scala 251:68]
  wire  _GEN_367; // @[TLB.scala 251:68]
  wire  _GEN_371; // @[TLB.scala 251:68]
  wire  _GEN_373; // @[TLB.scala 251:68]
  wire  _GEN_374; // @[TLB.scala 251:68]
  wire  _GEN_375; // @[TLB.scala 251:68]
  wire  _GEN_376; // @[TLB.scala 251:68]
  wire  _GEN_383; // @[TLB.scala 251:68]
  wire  _GEN_384; // @[TLB.scala 251:68]
  wire  _GEN_385; // @[TLB.scala 251:68]
  wire  _GEN_386; // @[TLB.scala 251:68]
  wire  _GEN_393; // @[TLB.scala 251:68]
  wire  _GEN_394; // @[TLB.scala 251:68]
  wire  _GEN_395; // @[TLB.scala 251:68]
  wire  _GEN_396; // @[TLB.scala 251:68]
  wire  _GEN_403; // @[TLB.scala 251:68]
  wire  _GEN_404; // @[TLB.scala 251:68]
  wire  _GEN_405; // @[TLB.scala 251:68]
  wire  _GEN_406; // @[TLB.scala 251:68]
  wire  _GEN_413; // @[TLB.scala 251:68]
  wire  _GEN_414; // @[TLB.scala 251:68]
  wire  _GEN_415; // @[TLB.scala 251:68]
  wire  _GEN_416; // @[TLB.scala 251:68]
  wire  _GEN_423; // @[TLB.scala 251:68]
  wire  _GEN_424; // @[TLB.scala 251:68]
  wire  _GEN_425; // @[TLB.scala 251:68]
  wire  _GEN_426; // @[TLB.scala 251:68]
  wire  _GEN_433; // @[TLB.scala 251:68]
  wire  _GEN_434; // @[TLB.scala 251:68]
  wire  _GEN_435; // @[TLB.scala 251:68]
  wire  _GEN_436; // @[TLB.scala 251:68]
  wire  _GEN_443; // @[TLB.scala 251:68]
  wire  _GEN_444; // @[TLB.scala 251:68]
  wire  _GEN_445; // @[TLB.scala 251:68]
  wire  _GEN_446; // @[TLB.scala 251:68]
  wire  _GEN_455; // @[TLB.scala 224:40]
  wire  _GEN_459; // @[TLB.scala 224:40]
  wire  _GEN_463; // @[TLB.scala 224:40]
  wire  _GEN_467; // @[TLB.scala 224:40]
  wire  _GEN_471; // @[TLB.scala 224:40]
  wire  _GEN_473; // @[TLB.scala 224:40]
  wire  _GEN_474; // @[TLB.scala 224:40]
  wire  _GEN_475; // @[TLB.scala 224:40]
  wire  _GEN_476; // @[TLB.scala 224:40]
  wire  _GEN_483; // @[TLB.scala 224:40]
  wire  _GEN_484; // @[TLB.scala 224:40]
  wire  _GEN_485; // @[TLB.scala 224:40]
  wire  _GEN_486; // @[TLB.scala 224:40]
  wire  _GEN_493; // @[TLB.scala 224:40]
  wire  _GEN_494; // @[TLB.scala 224:40]
  wire  _GEN_495; // @[TLB.scala 224:40]
  wire  _GEN_496; // @[TLB.scala 224:40]
  wire  _GEN_503; // @[TLB.scala 224:40]
  wire  _GEN_504; // @[TLB.scala 224:40]
  wire  _GEN_505; // @[TLB.scala 224:40]
  wire  _GEN_506; // @[TLB.scala 224:40]
  wire  _GEN_513; // @[TLB.scala 224:40]
  wire  _GEN_514; // @[TLB.scala 224:40]
  wire  _GEN_515; // @[TLB.scala 224:40]
  wire  _GEN_516; // @[TLB.scala 224:40]
  wire  _GEN_523; // @[TLB.scala 224:40]
  wire  _GEN_524; // @[TLB.scala 224:40]
  wire  _GEN_525; // @[TLB.scala 224:40]
  wire  _GEN_526; // @[TLB.scala 224:40]
  wire  _GEN_533; // @[TLB.scala 224:40]
  wire  _GEN_534; // @[TLB.scala 224:40]
  wire  _GEN_535; // @[TLB.scala 224:40]
  wire  _GEN_536; // @[TLB.scala 224:40]
  wire  _GEN_543; // @[TLB.scala 224:40]
  wire  _GEN_544; // @[TLB.scala 224:40]
  wire  _GEN_545; // @[TLB.scala 224:40]
  wire  _GEN_546; // @[TLB.scala 224:40]
  wire [5:0] _T_2136; // @[Cat.scala 30:58]
  wire [13:0] ptw_ae_array; // @[Cat.scala 30:58]
  wire  _T_2145; // @[TLB.scala 306:32]
  wire [5:0] _T_2150; // @[Cat.scala 30:58]
  wire [12:0] _T_2157; // @[Cat.scala 30:58]
  wire [12:0] _T_2158; // @[TLB.scala 306:23]
  wire [12:0] _T_2172; // @[TLB.scala 306:89]
  wire [12:0] priv_rw_ok; // @[TLB.scala 306:84]
  wire [5:0] _T_2202; // @[Cat.scala 30:58]
  wire [12:0] _T_2209; // @[Cat.scala 30:58]
  wire [5:0] _T_2214; // @[Cat.scala 30:58]
  wire [12:0] _T_2221; // @[Cat.scala 30:58]
  wire [12:0] _T_2222; // @[TLB.scala 308:73]
  wire [12:0] _T_2223; // @[TLB.scala 308:68]
  wire [12:0] _T_2224; // @[TLB.scala 308:40]
  wire [13:0] r_array; // @[Cat.scala 30:58]
  wire [5:0] _T_2229; // @[Cat.scala 30:58]
  wire [12:0] _T_2236; // @[Cat.scala 30:58]
  wire [12:0] _T_2237; // @[TLB.scala 309:40]
  wire [13:0] w_array; // @[Cat.scala 30:58]
  wire [1:0] _T_2252; // @[Bitwise.scala 72:12]
  wire [5:0] _T_2257; // @[Cat.scala 30:58]
  wire [13:0] _T_2264; // @[Cat.scala 30:58]
  wire [13:0] pr_array; // @[TLB.scala 311:87]
  wire [1:0] _T_2266; // @[Bitwise.scala 72:12]
  wire [5:0] _T_2271; // @[Cat.scala 30:58]
  wire [13:0] _T_2278; // @[Cat.scala 30:58]
  wire [13:0] pw_array; // @[TLB.scala 312:87]
  wire [1:0] _T_2294; // @[Bitwise.scala 72:12]
  wire [5:0] _T_2299; // @[Cat.scala 30:58]
  wire [13:0] paa_array; // @[Cat.scala 30:58]
  wire [5:0] _T_2312; // @[Cat.scala 30:58]
  wire [13:0] pal_array; // @[Cat.scala 30:58]
  wire [1:0] _T_2320; // @[Bitwise.scala 72:12]
  wire [5:0] _T_2325; // @[Cat.scala 30:58]
  wire [13:0] eff_array; // @[Cat.scala 30:58]
  wire [1:0] _T_2333; // @[Bitwise.scala 72:12]
  wire [5:0] _T_2338; // @[Cat.scala 30:58]
  wire [13:0] c_array; // @[Cat.scala 30:58]
  wire [3:0] _T_2358; // @[OneHot.scala 45:35]
  wire [3:0] _T_2361; // @[TLB.scala 320:69]
  wire [39:0] _GEN_1000; // @[TLB.scala 320:39]
  wire [39:0] _T_2362; // @[TLB.scala 320:39]
  wire  misaligned; // @[TLB.scala 320:75]
  wire  _T_2364; // @[TLB.scala 323:37]
  wire [26:0] _T_2365; // @[TLB.scala 323:53]
  wire  _T_2366; // @[TLB.scala 323:60]
  wire  _T_2367; // @[TLB.scala 323:44]
  wire  bad_va; // @[TLB.scala 321:27]
  wire [13:0] _T_2368; // @[TLB.scala 327:8]
  wire  _T_2369; // @[package.scala 14:47]
  wire  _T_2370; // @[package.scala 14:47]
  wire  _T_2371; // @[package.scala 14:62]
  wire [13:0] _T_2374; // @[TLB.scala 328:8]
  wire [13:0] ae_array; // @[TLB.scala 327:37]
  wire  _T_2375; // @[Consts.scala 93:31]
  wire  _T_2377; // @[Consts.scala 93:41]
  wire  _T_2379; // @[Consts.scala 93:58]
  wire  _T_2380; // @[package.scala 14:47]
  wire  _T_2381; // @[package.scala 14:47]
  wire  _T_2382; // @[package.scala 14:47]
  wire  _T_2383; // @[package.scala 14:47]
  wire  _T_2384; // @[package.scala 14:62]
  wire  _T_2385; // @[package.scala 14:62]
  wire  _T_2386; // @[package.scala 14:62]
  wire  _T_2387; // @[package.scala 14:47]
  wire  _T_2388; // @[package.scala 14:47]
  wire  _T_2389; // @[package.scala 14:47]
  wire  _T_2390; // @[package.scala 14:47]
  wire  _T_2391; // @[package.scala 14:47]
  wire  _T_2392; // @[package.scala 14:62]
  wire  _T_2393; // @[package.scala 14:62]
  wire  _T_2394; // @[package.scala 14:62]
  wire  _T_2395; // @[package.scala 14:62]
  wire  _T_2396; // @[Consts.scala 91:44]
  wire  _T_2397; // @[Consts.scala 93:75]
  wire [13:0] _T_2399; // @[TLB.scala 329:59]
  wire [13:0] ae_ld_array; // @[TLB.scala 329:24]
  wire  _T_2400; // @[Consts.scala 94:32]
  wire  _T_2401; // @[Consts.scala 94:49]
  wire  _T_2402; // @[Consts.scala 94:42]
  wire  _T_2404; // @[Consts.scala 94:59]
  wire  _T_2422; // @[Consts.scala 94:76]
  wire [13:0] _T_2424; // @[TLB.scala 331:44]
  wire [13:0] _T_2425; // @[TLB.scala 331:8]
  wire [13:0] _T_2435; // @[TLB.scala 332:8]
  wire [13:0] _T_2436; // @[TLB.scala 331:62]
  wire [13:0] _T_2448; // @[TLB.scala 333:8]
  wire [13:0] ae_st_array; // @[TLB.scala 332:79]
  wire  _T_2472; // @[TLB.scala 334:36]
  wire [13:0] ma_ld_array; // @[TLB.scala 334:24]
  wire  _T_2497; // @[TLB.scala 335:36]
  wire [13:0] ma_st_array; // @[TLB.scala 335:24]
  wire [13:0] _T_2522; // @[TLB.scala 336:60]
  wire [13:0] pf_ld_array; // @[TLB.scala 336:24]
  wire [13:0] _T_2547; // @[TLB.scala 337:61]
  wire [13:0] pf_st_array; // @[TLB.scala 337:24]
  wire  tlb_hit; // @[TLB.scala 340:27]
  wire  _T_2551; // @[TLB.scala 341:29]
  wire  tlb_miss; // @[TLB.scala 341:40]
  reg [6:0] _T_2554; // @[Replacement.scala 41:30]
  reg [31:0] _RAND_100;
  reg [2:0] _T_2556; // @[Replacement.scala 41:30]
  reg [31:0] _RAND_101;
  wire  _T_2557; // @[TLB.scala 345:22]
  wire  _T_2558; // @[package.scala 63:59]
  wire  _T_2559; // @[package.scala 63:59]
  wire  _T_2560; // @[package.scala 63:59]
  wire  _T_2561; // @[package.scala 63:59]
  wire  _T_2562; // @[package.scala 63:59]
  wire  _T_2563; // @[package.scala 63:59]
  wire  _T_2564; // @[package.scala 63:59]
  wire [7:0] _T_2571; // @[Cat.scala 30:58]
  wire  _T_2574; // @[OneHot.scala 28:14]
  wire [3:0] _T_2575; // @[OneHot.scala 28:28]
  wire  _T_2578; // @[OneHot.scala 28:14]
  wire [1:0] _T_2579; // @[OneHot.scala 28:28]
  wire [2:0] _T_2582; // @[Cat.scala 30:58]
  wire [7:0] _T_2583; // @[Replacement.scala 46:28]
  wire [7:0] _T_2587; // @[Replacement.scala 50:37]
  wire [7:0] _T_2589; // @[Replacement.scala 50:37]
  wire [7:0] _T_2591; // @[Replacement.scala 50:37]
  wire [1:0] _T_2592; // @[Cat.scala 30:58]
  wire [3:0] _T_2595; // @[Replacement.scala 50:37]
  wire [7:0] _GEN_1001; // @[Replacement.scala 50:37]
  wire [7:0] _T_2596; // @[Replacement.scala 50:37]
  wire [7:0] _T_2598; // @[Replacement.scala 50:37]
  wire [7:0] _T_2600; // @[Replacement.scala 50:37]
  wire [2:0] _T_2601; // @[Cat.scala 30:58]
  wire [7:0] _T_2604; // @[Replacement.scala 50:37]
  wire [7:0] _T_2605; // @[Replacement.scala 50:37]
  wire [7:0] _T_2607; // @[Replacement.scala 50:37]
  wire [7:0] _T_2609; // @[Replacement.scala 50:37]
  wire  _T_2612; // @[package.scala 63:59]
  wire  _T_2613; // @[package.scala 63:59]
  wire  _T_2614; // @[package.scala 63:59]
  wire [3:0] _T_2617; // @[Cat.scala 30:58]
  wire  _T_2620; // @[OneHot.scala 28:14]
  wire [1:0] _T_2621; // @[OneHot.scala 28:28]
  wire [1:0] _T_2623; // @[Cat.scala 30:58]
  wire [3:0] _T_2624; // @[Replacement.scala 46:28]
  wire [3:0] _T_2628; // @[Replacement.scala 50:37]
  wire [3:0] _T_2630; // @[Replacement.scala 50:37]
  wire [3:0] _T_2632; // @[Replacement.scala 50:37]
  wire [1:0] _T_2633; // @[Cat.scala 30:58]
  wire [3:0] _T_2636; // @[Replacement.scala 50:37]
  wire [3:0] _T_2637; // @[Replacement.scala 50:37]
  wire [3:0] _T_2639; // @[Replacement.scala 50:37]
  wire [3:0] _T_2641; // @[Replacement.scala 50:37]
  wire  _T_2653; // @[Misc.scala 187:16]
  wire  _T_2655; // @[Misc.scala 187:61]
  wire  _T_2657; // @[Misc.scala 187:16]
  wire  _T_2659; // @[Misc.scala 187:61]
  wire  _T_2660; // @[Misc.scala 187:49]
  wire  _T_2669; // @[Misc.scala 187:16]
  wire  _T_2671; // @[Misc.scala 187:61]
  wire  _T_2673; // @[Misc.scala 187:16]
  wire  _T_2675; // @[Misc.scala 187:61]
  wire  _T_2676; // @[Misc.scala 187:49]
  wire  _T_2677; // @[Misc.scala 187:16]
  wire  _T_2678; // @[Misc.scala 187:37]
  wire  _T_2679; // @[Misc.scala 187:61]
  wire  _T_2680; // @[Misc.scala 187:49]
  wire  _T_2690; // @[Misc.scala 187:16]
  wire  _T_2692; // @[Misc.scala 187:61]
  wire  _T_2694; // @[Misc.scala 187:16]
  wire  _T_2696; // @[Misc.scala 187:61]
  wire  _T_2697; // @[Misc.scala 187:49]
  wire  _T_2704; // @[Misc.scala 187:16]
  wire  _T_2706; // @[Misc.scala 187:61]
  wire  _T_2713; // @[Misc.scala 187:16]
  wire  _T_2715; // @[Misc.scala 187:61]
  wire  _T_2717; // @[Misc.scala 187:16]
  wire  _T_2718; // @[Misc.scala 187:37]
  wire  _T_2719; // @[Misc.scala 187:61]
  wire  _T_2720; // @[Misc.scala 187:49]
  wire  _T_2721; // @[Misc.scala 187:16]
  wire  _T_2722; // @[Misc.scala 187:37]
  wire  _T_2723; // @[Misc.scala 187:61]
  wire  _T_2724; // @[Misc.scala 187:49]
  wire  _T_2726; // @[Misc.scala 187:37]
  wire  _T_2727; // @[Misc.scala 187:61]
  wire  multipleHits; // @[Misc.scala 187:49]
  wire  _T_2752; // @[TLB.scala 358:28]
  wire [13:0] _T_2753; // @[TLB.scala 358:72]
  wire  _T_2754; // @[TLB.scala 358:80]
  wire  _T_2779; // @[TLB.scala 359:28]
  wire [13:0] _T_2780; // @[TLB.scala 359:73]
  wire  _T_2781; // @[TLB.scala 359:81]
  wire [13:0] _T_2786; // @[TLB.scala 361:33]
  wire [13:0] _T_2788; // @[TLB.scala 362:33]
  wire [13:0] _T_2793; // @[TLB.scala 364:33]
  wire [13:0] _T_2795; // @[TLB.scala 365:33]
  wire [13:0] _T_2797; // @[TLB.scala 367:33]
  wire  _T_2802; // @[TLB.scala 369:29]
  wire  _T_2808; // @[Decoupled.scala 37:37]
  wire  _T_2809; // @[TLB.scala 385:25]
  wire [3:0] _T_2814; // @[Replacement.scala 61:48]
  wire [1:0] _T_2817; // @[Cat.scala 30:58]
  wire [3:0] _T_2821; // @[Replacement.scala 61:48]
  wire [2:0] _T_2824; // @[Cat.scala 30:58]
  wire [3:0] _T_2828; // @[Cat.scala 30:58]
  wire  _T_2830; // @[TLB.scala 440:16]
  wire  _T_2832; // @[OneHot.scala 39:40]
  wire  _T_2833; // @[OneHot.scala 39:40]
  wire  _T_2834; // @[OneHot.scala 39:40]
  wire [7:0] _T_2844; // @[Replacement.scala 61:48]
  wire [1:0] _T_2847; // @[Cat.scala 30:58]
  wire [7:0] _T_2851; // @[Replacement.scala 61:48]
  wire [2:0] _T_2854; // @[Cat.scala 30:58]
  wire [7:0] _T_2858; // @[Replacement.scala 61:48]
  wire [3:0] _T_2861; // @[Cat.scala 30:58]
  wire [7:0] _T_2893; // @[Cat.scala 30:58]
  wire  _T_2895; // @[TLB.scala 440:16]
  wire  _T_2897; // @[OneHot.scala 39:40]
  wire  _T_2898; // @[OneHot.scala 39:40]
  wire  _T_2899; // @[OneHot.scala 39:40]
  wire  _T_2900; // @[OneHot.scala 39:40]
  wire  _T_2901; // @[OneHot.scala 39:40]
  wire  _T_2902; // @[OneHot.scala 39:40]
  wire  _T_2903; // @[OneHot.scala 39:40]
  wire  _T_2940; // @[TLB.scala 399:17]
  wire  _T_2941; // @[TLB.scala 399:28]
  wire  _T_2946; // @[TLB.scala 414:72]
  wire  _T_2947; // @[TLB.scala 414:34]
  wire  _T_2949; // @[TLB.scala 414:13]
  wire  _T_2957; // @[TLB.scala 150:63]
  wire  _GEN_652; // @[TLB.scala 158:21]
  wire  _GEN_653; // @[TLB.scala 158:21]
  wire  _GEN_654; // @[TLB.scala 158:21]
  wire  _GEN_655; // @[TLB.scala 158:21]
  wire  _GEN_656; // @[TLB.scala 417:40]
  wire  _GEN_657; // @[TLB.scala 417:40]
  wire  _GEN_658; // @[TLB.scala 417:40]
  wire  _GEN_659; // @[TLB.scala 417:40]
  wire  _T_3128; // @[TLB.scala 150:63]
  wire  _GEN_680; // @[TLB.scala 158:21]
  wire  _GEN_681; // @[TLB.scala 158:21]
  wire  _GEN_682; // @[TLB.scala 158:21]
  wire  _GEN_683; // @[TLB.scala 158:21]
  wire  _GEN_684; // @[TLB.scala 417:40]
  wire  _GEN_685; // @[TLB.scala 417:40]
  wire  _GEN_686; // @[TLB.scala 417:40]
  wire  _GEN_687; // @[TLB.scala 417:40]
  wire  _T_3299; // @[TLB.scala 150:63]
  wire  _GEN_708; // @[TLB.scala 158:21]
  wire  _GEN_709; // @[TLB.scala 158:21]
  wire  _GEN_710; // @[TLB.scala 158:21]
  wire  _GEN_711; // @[TLB.scala 158:21]
  wire  _GEN_712; // @[TLB.scala 417:40]
  wire  _GEN_713; // @[TLB.scala 417:40]
  wire  _GEN_714; // @[TLB.scala 417:40]
  wire  _GEN_715; // @[TLB.scala 417:40]
  wire  _T_3470; // @[TLB.scala 150:63]
  wire  _GEN_736; // @[TLB.scala 158:21]
  wire  _GEN_737; // @[TLB.scala 158:21]
  wire  _GEN_738; // @[TLB.scala 158:21]
  wire  _GEN_739; // @[TLB.scala 158:21]
  wire  _GEN_740; // @[TLB.scala 417:40]
  wire  _GEN_741; // @[TLB.scala 417:40]
  wire  _GEN_742; // @[TLB.scala 417:40]
  wire  _GEN_743; // @[TLB.scala 417:40]
  wire  _T_3641; // @[TLB.scala 150:63]
  wire  _GEN_764; // @[TLB.scala 158:21]
  wire  _GEN_765; // @[TLB.scala 158:21]
  wire  _GEN_766; // @[TLB.scala 158:21]
  wire  _GEN_767; // @[TLB.scala 158:21]
  wire  _GEN_768; // @[TLB.scala 417:40]
  wire  _GEN_769; // @[TLB.scala 417:40]
  wire  _GEN_770; // @[TLB.scala 417:40]
  wire  _GEN_771; // @[TLB.scala 417:40]
  wire  _T_3812; // @[TLB.scala 150:63]
  wire  _GEN_792; // @[TLB.scala 158:21]
  wire  _GEN_793; // @[TLB.scala 158:21]
  wire  _GEN_794; // @[TLB.scala 158:21]
  wire  _GEN_795; // @[TLB.scala 158:21]
  wire  _GEN_796; // @[TLB.scala 417:40]
  wire  _GEN_797; // @[TLB.scala 417:40]
  wire  _GEN_798; // @[TLB.scala 417:40]
  wire  _GEN_799; // @[TLB.scala 417:40]
  wire  _T_3983; // @[TLB.scala 150:63]
  wire  _GEN_820; // @[TLB.scala 158:21]
  wire  _GEN_821; // @[TLB.scala 158:21]
  wire  _GEN_822; // @[TLB.scala 158:21]
  wire  _GEN_823; // @[TLB.scala 158:21]
  wire  _GEN_824; // @[TLB.scala 417:40]
  wire  _GEN_825; // @[TLB.scala 417:40]
  wire  _GEN_826; // @[TLB.scala 417:40]
  wire  _GEN_827; // @[TLB.scala 417:40]
  wire  _T_4154; // @[TLB.scala 150:63]
  wire  _GEN_848; // @[TLB.scala 158:21]
  wire  _GEN_849; // @[TLB.scala 158:21]
  wire  _GEN_850; // @[TLB.scala 158:21]
  wire  _GEN_851; // @[TLB.scala 158:21]
  wire  _GEN_852; // @[TLB.scala 417:40]
  wire  _GEN_853; // @[TLB.scala 417:40]
  wire  _GEN_854; // @[TLB.scala 417:40]
  wire  _GEN_855; // @[TLB.scala 417:40]
  wire  _GEN_861; // @[TLB.scala 158:21]
  wire  _GEN_862; // @[TLB.scala 417:40]
  wire  _GEN_865; // @[TLB.scala 158:21]
  wire  _GEN_866; // @[TLB.scala 417:40]
  wire  _GEN_869; // @[TLB.scala 158:21]
  wire  _GEN_870; // @[TLB.scala 417:40]
  wire  _GEN_873; // @[TLB.scala 158:21]
  wire  _GEN_874; // @[TLB.scala 417:40]
  wire  _GEN_877; // @[TLB.scala 158:21]
  wire  _GEN_878; // @[TLB.scala 417:40]
  wire  _T_4530; // @[TLB.scala 421:24]
  reg [19:0] TLB_state; // @[Register tracking TLB state]
  reg [31:0] _RAND_102;
  reg  TLB_cov [0:1048575]; // @[Coverage map for TLB]
  reg [31:0] _RAND_103;
  wire  TLB_cov_read_data; // @[Coverage map for TLB]
  wire [19:0] TLB_cov_read_addr; // @[Coverage map for TLB]
  wire  TLB_cov_write_data; // @[Coverage map for TLB]
  wire [19:0] TLB_cov_write_addr; // @[Coverage map for TLB]
  wire  TLB_cov_write_mask; // @[Coverage map for TLB]
  wire  TLB_cov_write_en; // @[Coverage map for TLB]
  reg [29:0] TLB_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_104;
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  mux_cond_4;
  wire  mux_cond_5;
  wire  mux_cond_6;
  wire  mux_cond_7;
  wire  mux_cond_8;
  wire  mux_cond_9;
  wire  mux_cond_10;
  wire  mux_cond_11;
  wire  mux_cond_12;
  wire  mux_cond_13;
  wire  mux_cond_14;
  wire  mux_cond_15;
  wire  mux_cond_16;
  wire  mux_cond_17;
  wire  mux_cond_18;
  wire  mux_cond_19;
  wire  mux_cond_20;
  wire  mux_cond_21;
  wire  mux_cond_22;
  wire  mux_cond_23;
  wire  mux_cond_24;
  wire  mux_cond_25;
  wire  mux_cond_26;
  wire  mux_cond_27;
  wire  mux_cond_28;
  wire  mux_cond_29;
  wire  mux_cond_30;
  wire  mux_cond_31;
  wire  mux_cond_32;
  wire  mux_cond_33;
  wire  mux_cond_34;
  wire  mux_cond_35;
  wire  mux_cond_36;
  wire  mux_cond_37;
  wire  mux_cond_38;
  wire  mux_cond_39;
  wire  mux_cond_40;
  wire  mux_cond_41;
  wire  mux_cond_42;
  wire  mux_cond_43;
  wire  mux_cond_44;
  wire  mux_cond_45;
  wire  mux_cond_46;
  wire  mux_cond_47;
  wire  mux_cond_48;
  wire  mux_cond_49;
  wire  mux_cond_50;
  wire  mux_cond_51;
  wire  mux_cond_52;
  wire  mux_cond_53;
  wire  mux_cond_54;
  wire  mux_cond_55;
  wire  mux_cond_56;
  wire  mux_cond_57;
  wire  mux_cond_58;
  wire  mux_cond_59;
  wire  mux_cond_60;
  wire  mux_cond_61;
  wire  mux_cond_62;
  wire  mux_cond_63;
  wire  mux_cond_64;
  wire  mux_cond_65;
  wire  mux_cond_66;
  wire  mux_cond_67;
  wire  mux_cond_68;
  wire  mux_cond_69;
  wire  mux_cond_70;
  wire  mux_cond_71;
  wire  mux_cond_72;
  wire  mux_cond_73;
  wire [9:0] r_superpage_repl_addr_shl;
  wire [19:0] r_superpage_repl_addr_pad;
  wire [2:0] state_shl;
  wire [19:0] state_pad;
  wire [15:0] r_sectored_repl_addr_shl;
  wire [19:0] r_sectored_repl_addr_pad;
  wire [7:0] r_sectored_hit_addr_shl;
  wire [19:0] r_sectored_hit_addr_pad;
  wire [10:0] special_entry_valid_0_shl;
  wire [19:0] special_entry_valid_0_pad;
  wire [1:0] special_entry_level_shl;
  wire [19:0] special_entry_level_pad;
  wire [19:0] r_sectored_hit_shl;
  wire [19:0] r_sectored_hit_pad;
  wire [9:0] mux_cond_0_shl;
  wire [19:0] mux_cond_0_pad;
  wire [18:0] mux_cond_1_shl;
  wire [19:0] mux_cond_1_pad;
  wire [4:0] mux_cond_2_shl;
  wire [19:0] mux_cond_2_pad;
  wire [5:0] mux_cond_3_shl;
  wire [19:0] mux_cond_3_pad;
  wire [15:0] mux_cond_4_shl;
  wire [19:0] mux_cond_4_pad;
  wire [2:0] mux_cond_5_shl;
  wire [19:0] mux_cond_5_pad;
  wire [1:0] mux_cond_6_shl;
  wire [19:0] mux_cond_6_pad;
  wire [9:0] mux_cond_7_shl;
  wire [19:0] mux_cond_7_pad;
  wire [5:0] mux_cond_8_shl;
  wire [19:0] mux_cond_8_pad;
  wire [5:0] mux_cond_9_shl;
  wire [19:0] mux_cond_9_pad;
  wire [7:0] mux_cond_10_shl;
  wire [19:0] mux_cond_10_pad;
  wire [1:0] mux_cond_11_shl;
  wire [19:0] mux_cond_11_pad;
  wire [14:0] mux_cond_12_shl;
  wire [19:0] mux_cond_12_pad;
  wire [11:0] mux_cond_13_shl;
  wire [19:0] mux_cond_13_pad;
  wire [2:0] mux_cond_14_shl;
  wire [19:0] mux_cond_14_pad;
  wire [17:0] mux_cond_15_shl;
  wire [19:0] mux_cond_15_pad;
  wire  mux_cond_16_shl;
  wire [19:0] mux_cond_16_pad;
  wire [18:0] mux_cond_17_shl;
  wire [19:0] mux_cond_17_pad;
  wire [19:0] mux_cond_18_shl;
  wire [19:0] mux_cond_18_pad;
  wire [8:0] mux_cond_19_shl;
  wire [19:0] mux_cond_19_pad;
  wire [17:0] mux_cond_20_shl;
  wire [19:0] mux_cond_20_pad;
  wire [3:0] mux_cond_21_shl;
  wire [19:0] mux_cond_21_pad;
  wire [5:0] mux_cond_22_shl;
  wire [19:0] mux_cond_22_pad;
  wire [5:0] mux_cond_23_shl;
  wire [19:0] mux_cond_23_pad;
  wire [15:0] mux_cond_24_shl;
  wire [19:0] mux_cond_24_pad;
  wire [18:0] mux_cond_25_shl;
  wire [19:0] mux_cond_25_pad;
  wire [3:0] mux_cond_26_shl;
  wire [19:0] mux_cond_26_pad;
  wire [12:0] mux_cond_27_shl;
  wire [19:0] mux_cond_27_pad;
  wire [10:0] mux_cond_28_shl;
  wire [19:0] mux_cond_28_pad;
  wire [3:0] mux_cond_29_shl;
  wire [19:0] mux_cond_29_pad;
  wire  mux_cond_30_shl;
  wire [19:0] mux_cond_30_pad;
  wire [18:0] mux_cond_31_shl;
  wire [19:0] mux_cond_31_pad;
  wire [12:0] mux_cond_32_shl;
  wire [19:0] mux_cond_32_pad;
  wire [1:0] mux_cond_33_shl;
  wire [19:0] mux_cond_33_pad;
  wire [1:0] mux_cond_34_shl;
  wire [19:0] mux_cond_34_pad;
  wire [3:0] mux_cond_35_shl;
  wire [19:0] mux_cond_35_pad;
  wire [7:0] mux_cond_36_shl;
  wire [19:0] mux_cond_36_pad;
  wire [6:0] mux_cond_37_shl;
  wire [19:0] mux_cond_37_pad;
  wire [5:0] mux_cond_38_shl;
  wire [19:0] mux_cond_38_pad;
  wire [4:0] mux_cond_39_shl;
  wire [19:0] mux_cond_39_pad;
  wire [3:0] mux_cond_40_shl;
  wire [19:0] mux_cond_40_pad;
  wire [10:0] mux_cond_41_shl;
  wire [19:0] mux_cond_41_pad;
  wire [14:0] mux_cond_42_shl;
  wire [19:0] mux_cond_42_pad;
  wire [16:0] mux_cond_43_shl;
  wire [19:0] mux_cond_43_pad;
  wire [2:0] mux_cond_44_shl;
  wire [19:0] mux_cond_44_pad;
  wire [13:0] mux_cond_45_shl;
  wire [19:0] mux_cond_45_pad;
  wire [4:0] mux_cond_46_shl;
  wire [19:0] mux_cond_46_pad;
  wire [8:0] mux_cond_47_shl;
  wire [19:0] mux_cond_47_pad;
  wire [10:0] mux_cond_48_shl;
  wire [19:0] mux_cond_48_pad;
  wire [8:0] mux_cond_49_shl;
  wire [19:0] mux_cond_49_pad;
  wire [16:0] mux_cond_50_shl;
  wire [19:0] mux_cond_50_pad;
  wire [12:0] mux_cond_51_shl;
  wire [19:0] mux_cond_51_pad;
  wire [19:0] mux_cond_52_shl;
  wire [19:0] mux_cond_52_pad;
  wire [16:0] mux_cond_53_shl;
  wire [19:0] mux_cond_53_pad;
  wire [19:0] mux_cond_54_shl;
  wire [19:0] mux_cond_54_pad;
  wire [10:0] mux_cond_55_shl;
  wire [19:0] mux_cond_55_pad;
  wire [7:0] mux_cond_56_shl;
  wire [19:0] mux_cond_56_pad;
  wire [1:0] mux_cond_57_shl;
  wire [19:0] mux_cond_57_pad;
  wire [13:0] mux_cond_58_shl;
  wire [19:0] mux_cond_58_pad;
  wire [18:0] mux_cond_59_shl;
  wire [19:0] mux_cond_59_pad;
  wire [14:0] mux_cond_60_shl;
  wire [19:0] mux_cond_60_pad;
  wire [2:0] mux_cond_61_shl;
  wire [19:0] mux_cond_61_pad;
  wire [17:0] mux_cond_62_shl;
  wire [19:0] mux_cond_62_pad;
  wire [3:0] mux_cond_63_shl;
  wire [19:0] mux_cond_63_pad;
  wire [14:0] mux_cond_64_shl;
  wire [19:0] mux_cond_64_pad;
  wire [7:0] mux_cond_65_shl;
  wire [19:0] mux_cond_65_pad;
  wire [15:0] mux_cond_66_shl;
  wire [19:0] mux_cond_66_pad;
  wire [16:0] mux_cond_67_shl;
  wire [19:0] mux_cond_67_pad;
  wire [12:0] mux_cond_68_shl;
  wire [19:0] mux_cond_68_pad;
  wire [1:0] mux_cond_69_shl;
  wire [19:0] mux_cond_69_pad;
  wire [5:0] mux_cond_70_shl;
  wire [19:0] mux_cond_70_pad;
  wire [11:0] mux_cond_71_shl;
  wire [19:0] mux_cond_71_pad;
  wire [13:0] mux_cond_72_shl;
  wire [19:0] mux_cond_72_pad;
  wire [13:0] mux_cond_73_shl;
  wire [19:0] mux_cond_73_pad;
  wire [2:0] sectored_entries_7_valid_1_shl;
  wire [19:0] sectored_entries_7_valid_1_pad;
  wire [13:0] sectored_entries_5_valid_3_shl;
  wire [19:0] sectored_entries_5_valid_3_pad;
  wire [2:0] sectored_entries_5_valid_1_shl;
  wire [19:0] sectored_entries_5_valid_1_pad;
  wire [2:0] sectored_entries_4_valid_1_shl;
  wire [19:0] sectored_entries_4_valid_1_pad;
  wire [5:0] superpage_entries_0_valid_0_shl;
  wire [19:0] superpage_entries_0_valid_0_pad;
  wire [17:0] sectored_entries_3_valid_2_shl;
  wire [19:0] sectored_entries_3_valid_2_pad;
  wire [17:0] sectored_entries_1_valid_0_shl;
  wire [19:0] sectored_entries_1_valid_0_pad;
  wire [11:0] superpage_entries_3_level_shl;
  wire [19:0] superpage_entries_3_level_pad;
  wire [17:0] sectored_entries_5_valid_0_shl;
  wire [19:0] sectored_entries_5_valid_0_pad;
  wire [2:0] sectored_entries_0_valid_1_shl;
  wire [19:0] sectored_entries_0_valid_1_pad;
  wire [17:0] sectored_entries_3_valid_0_shl;
  wire [19:0] sectored_entries_3_valid_0_pad;
  wire [17:0] sectored_entries_7_valid_2_shl;
  wire [19:0] sectored_entries_7_valid_2_pad;
  wire [13:0] sectored_entries_2_valid_3_shl;
  wire [19:0] sectored_entries_2_valid_3_pad;
  wire [17:0] sectored_entries_4_valid_0_shl;
  wire [19:0] sectored_entries_4_valid_0_pad;
  wire [13:0] sectored_entries_6_valid_3_shl;
  wire [19:0] sectored_entries_6_valid_3_pad;
  wire [13:0] sectored_entries_1_valid_3_shl;
  wire [19:0] sectored_entries_1_valid_3_pad;
  wire [17:0] sectored_entries_6_valid_0_shl;
  wire [19:0] sectored_entries_6_valid_0_pad;
  wire [17:0] sectored_entries_2_valid_2_shl;
  wire [19:0] sectored_entries_2_valid_2_pad;
  wire [17:0] sectored_entries_6_valid_2_shl;
  wire [19:0] sectored_entries_6_valid_2_pad;
  wire [2:0] sectored_entries_6_valid_1_shl;
  wire [19:0] sectored_entries_6_valid_1_pad;
  wire [13:0] sectored_entries_4_valid_3_shl;
  wire [19:0] sectored_entries_4_valid_3_pad;
  wire [17:0] sectored_entries_1_valid_2_shl;
  wire [19:0] sectored_entries_1_valid_2_pad;
  wire [17:0] sectored_entries_5_valid_2_shl;
  wire [19:0] sectored_entries_5_valid_2_pad;
  wire [11:0] superpage_entries_2_level_shl;
  wire [19:0] superpage_entries_2_level_pad;
  wire [5:0] superpage_entries_3_valid_0_shl;
  wire [19:0] superpage_entries_3_valid_0_pad;
  wire [2:0] sectored_entries_1_valid_1_shl;
  wire [19:0] sectored_entries_1_valid_1_pad;
  wire [17:0] sectored_entries_0_valid_0_shl;
  wire [19:0] sectored_entries_0_valid_0_pad;
  wire [5:0] superpage_entries_1_valid_0_shl;
  wire [19:0] superpage_entries_1_valid_0_pad;
  wire [13:0] sectored_entries_0_valid_3_shl;
  wire [19:0] sectored_entries_0_valid_3_pad;
  wire [17:0] sectored_entries_7_valid_0_shl;
  wire [19:0] sectored_entries_7_valid_0_pad;
  wire [17:0] sectored_entries_0_valid_2_shl;
  wire [19:0] sectored_entries_0_valid_2_pad;
  wire [11:0] superpage_entries_0_level_shl;
  wire [19:0] superpage_entries_0_level_pad;
  wire [2:0] sectored_entries_2_valid_1_shl;
  wire [19:0] sectored_entries_2_valid_1_pad;
  wire [2:0] sectored_entries_3_valid_1_shl;
  wire [19:0] sectored_entries_3_valid_1_pad;
  wire [17:0] sectored_entries_2_valid_0_shl;
  wire [19:0] sectored_entries_2_valid_0_pad;
  wire [13:0] sectored_entries_7_valid_3_shl;
  wire [19:0] sectored_entries_7_valid_3_pad;
  wire [17:0] sectored_entries_4_valid_2_shl;
  wire [19:0] sectored_entries_4_valid_2_pad;
  wire [13:0] sectored_entries_3_valid_3_shl;
  wire [19:0] sectored_entries_3_valid_3_pad;
  wire [11:0] superpage_entries_1_level_shl;
  wire [19:0] superpage_entries_1_level_pad;
  wire [5:0] superpage_entries_2_valid_0_shl;
  wire [19:0] superpage_entries_2_valid_0_pad;
  wire [19:0] TLB_xor64;
  wire [19:0] TLB_xor31;
  wire [19:0] TLB_xor65;
  wire [19:0] TLB_xor66;
  wire [19:0] TLB_xor32;
  wire [19:0] TLB_xor15;
  wire [19:0] TLB_xor67;
  wire [19:0] TLB_xor68;
  wire [19:0] TLB_xor33;
  wire [19:0] TLB_xor69;
  wire [19:0] TLB_xor70;
  wire [19:0] TLB_xor34;
  wire [19:0] TLB_xor16;
  wire [19:0] TLB_xor7;
  wire [19:0] TLB_xor72;
  wire [19:0] TLB_xor35;
  wire [19:0] TLB_xor73;
  wire [19:0] TLB_xor74;
  wire [19:0] TLB_xor36;
  wire [19:0] TLB_xor17;
  wire [19:0] TLB_xor75;
  wire [19:0] TLB_xor76;
  wire [19:0] TLB_xor37;
  wire [19:0] TLB_xor77;
  wire [19:0] TLB_xor78;
  wire [19:0] TLB_xor38;
  wire [19:0] TLB_xor18;
  wire [19:0] TLB_xor8;
  wire [19:0] TLB_xor3;
  wire [19:0] TLB_xor80;
  wire [19:0] TLB_xor39;
  wire [19:0] TLB_xor81;
  wire [19:0] TLB_xor82;
  wire [19:0] TLB_xor40;
  wire [19:0] TLB_xor19;
  wire [19:0] TLB_xor83;
  wire [19:0] TLB_xor84;
  wire [19:0] TLB_xor41;
  wire [19:0] TLB_xor85;
  wire [19:0] TLB_xor86;
  wire [19:0] TLB_xor42;
  wire [19:0] TLB_xor20;
  wire [19:0] TLB_xor9;
  wire [19:0] TLB_xor88;
  wire [19:0] TLB_xor43;
  wire [19:0] TLB_xor89;
  wire [19:0] TLB_xor90;
  wire [19:0] TLB_xor44;
  wire [19:0] TLB_xor21;
  wire [19:0] TLB_xor91;
  wire [19:0] TLB_xor92;
  wire [19:0] TLB_xor45;
  wire [19:0] TLB_xor93;
  wire [19:0] TLB_xor94;
  wire [19:0] TLB_xor46;
  wire [19:0] TLB_xor22;
  wire [19:0] TLB_xor10;
  wire [19:0] TLB_xor4;
  wire [19:0] TLB_xor1;
  wire [19:0] TLB_xor96;
  wire [19:0] TLB_xor47;
  wire [19:0] TLB_xor97;
  wire [19:0] TLB_xor98;
  wire [19:0] TLB_xor48;
  wire [19:0] TLB_xor23;
  wire [19:0] TLB_xor99;
  wire [19:0] TLB_xor100;
  wire [19:0] TLB_xor49;
  wire [19:0] TLB_xor101;
  wire [19:0] TLB_xor102;
  wire [19:0] TLB_xor50;
  wire [19:0] TLB_xor24;
  wire [19:0] TLB_xor11;
  wire [19:0] TLB_xor104;
  wire [19:0] TLB_xor51;
  wire [19:0] TLB_xor105;
  wire [19:0] TLB_xor106;
  wire [19:0] TLB_xor52;
  wire [19:0] TLB_xor25;
  wire [19:0] TLB_xor107;
  wire [19:0] TLB_xor108;
  wire [19:0] TLB_xor53;
  wire [19:0] TLB_xor109;
  wire [19:0] TLB_xor110;
  wire [19:0] TLB_xor54;
  wire [19:0] TLB_xor26;
  wire [19:0] TLB_xor12;
  wire [19:0] TLB_xor5;
  wire [19:0] TLB_xor112;
  wire [19:0] TLB_xor55;
  wire [19:0] TLB_xor113;
  wire [19:0] TLB_xor114;
  wire [19:0] TLB_xor56;
  wire [19:0] TLB_xor27;
  wire [19:0] TLB_xor115;
  wire [19:0] TLB_xor116;
  wire [19:0] TLB_xor57;
  wire [19:0] TLB_xor117;
  wire [19:0] TLB_xor118;
  wire [19:0] TLB_xor58;
  wire [19:0] TLB_xor28;
  wire [19:0] TLB_xor13;
  wire [19:0] TLB_xor119;
  wire [19:0] TLB_xor120;
  wire [19:0] TLB_xor59;
  wire [19:0] TLB_xor121;
  wire [19:0] TLB_xor122;
  wire [19:0] TLB_xor60;
  wire [19:0] TLB_xor29;
  wire [19:0] TLB_xor123;
  wire [19:0] TLB_xor124;
  wire [19:0] TLB_xor61;
  wire [19:0] TLB_xor125;
  wire [19:0] TLB_xor126;
  wire [19:0] TLB_xor62;
  wire [19:0] TLB_xor30;
  wire [19:0] TLB_xor14;
  wire [19:0] TLB_xor6;
  wire [19:0] TLB_xor2;
  wire [19:0] TLB_xor0;
  wire [29:0] pmp_sum;
  wire  stopEn0;
  wire  pmp_metaAssert_wire;
  wire  TLB_or0;
  reg  TLB_metaAssert;
  reg [31:0] _RAND_105;
  PMPChecker pmp ( // @[TLB.scala 190:19]
    .io_prv(pmp_io_prv),
    .io_pmp_0_cfg_l(pmp_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(pmp_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(pmp_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(pmp_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(pmp_io_pmp_0_cfg_r),
    .io_pmp_0_addr(pmp_io_pmp_0_addr),
    .io_pmp_0_mask(pmp_io_pmp_0_mask),
    .io_pmp_1_cfg_l(pmp_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(pmp_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(pmp_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(pmp_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(pmp_io_pmp_1_cfg_r),
    .io_pmp_1_addr(pmp_io_pmp_1_addr),
    .io_pmp_1_mask(pmp_io_pmp_1_mask),
    .io_pmp_2_cfg_l(pmp_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(pmp_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(pmp_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(pmp_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(pmp_io_pmp_2_cfg_r),
    .io_pmp_2_addr(pmp_io_pmp_2_addr),
    .io_pmp_2_mask(pmp_io_pmp_2_mask),
    .io_pmp_3_cfg_l(pmp_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(pmp_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(pmp_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(pmp_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(pmp_io_pmp_3_cfg_r),
    .io_pmp_3_addr(pmp_io_pmp_3_addr),
    .io_pmp_3_mask(pmp_io_pmp_3_mask),
    .io_pmp_4_cfg_l(pmp_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(pmp_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(pmp_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(pmp_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(pmp_io_pmp_4_cfg_r),
    .io_pmp_4_addr(pmp_io_pmp_4_addr),
    .io_pmp_4_mask(pmp_io_pmp_4_mask),
    .io_pmp_5_cfg_l(pmp_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(pmp_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(pmp_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(pmp_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(pmp_io_pmp_5_cfg_r),
    .io_pmp_5_addr(pmp_io_pmp_5_addr),
    .io_pmp_5_mask(pmp_io_pmp_5_mask),
    .io_pmp_6_cfg_l(pmp_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(pmp_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(pmp_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(pmp_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(pmp_io_pmp_6_cfg_r),
    .io_pmp_6_addr(pmp_io_pmp_6_addr),
    .io_pmp_6_mask(pmp_io_pmp_6_mask),
    .io_pmp_7_cfg_l(pmp_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(pmp_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(pmp_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(pmp_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(pmp_io_pmp_7_cfg_r),
    .io_pmp_7_addr(pmp_io_pmp_7_addr),
    .io_pmp_7_mask(pmp_io_pmp_7_mask),
    .io_addr(pmp_io_addr),
    .io_size(pmp_io_size),
    .io_r(pmp_io_r),
    .io_w(pmp_io_w),
    .io_x(pmp_io_x),
    .io_covSum(pmp_io_covSum),
    .metaAssert(pmp_metaAssert)
  );
  assign priv_s = io_ptw_status_dprv[0]; // @[TLB.scala 178:20]
  assign priv_uses_vm = io_ptw_status_dprv <= 2'h1; // @[TLB.scala 179:27]
  assign _T_322 = io_ptw_ptbr_mode[3] & priv_uses_vm; // @[TLB.scala 180:83]
  assign vm_enabled = _T_322 & ~io_req_bits_passthrough; // @[TLB.scala 180:99]
  assign vpn = io_req_bits_vaddr[38:12]; // @[TLB.scala 183:30]
  assign refill_ppn = io_ptw_resp_bits_pte_ppn[19:0]; // @[TLB.scala 184:44]
  assign _T_324 = state == 2'h1; // @[package.scala 14:47]
  assign _T_325 = state == 2'h3; // @[package.scala 14:47]
  assign invalidate_refill = _T_324 | _T_325; // @[package.scala 14:62]
  assign _T_348 = special_entry_level < 2'h1; // @[TLB.scala 123:30]
  assign _T_350 = _T_348 ? vpn : 27'h0; // @[TLB.scala 124:30]
  assign _GEN_954 = {{7'd0}, special_entry_data_0[33:14]}; // @[TLB.scala 124:49]
  assign _T_351 = _T_350 | _GEN_954; // @[TLB.scala 124:49]
  assign _T_354 = special_entry_level < 2'h2; // @[TLB.scala 123:30]
  assign _T_356 = _T_354 ? vpn : 27'h0; // @[TLB.scala 124:30]
  assign _T_357 = _T_356 | _GEN_954; // @[TLB.scala 124:49]
  assign _T_359 = {special_entry_data_0[33:32],_T_351[17:9],_T_357[8:0]}; // @[Cat.scala 30:58]
  assign _T_361 = vm_enabled ? {{8'd0}, _T_359} : io_req_bits_vaddr[39:12]; // @[TLB.scala 188:20]
  assign mpu_ppn = io_ptw_resp_valid ? {{8'd0}, refill_ppn} : _T_361; // @[TLB.scala 187:20]
  assign mpu_physaddr = {mpu_ppn,io_req_bits_vaddr[11:0]}; // @[Cat.scala 30:58]
  assign _T_363 = io_ptw_resp_valid | io_req_bits_passthrough; // @[TLB.scala 194:49]
  assign _T_366 = mpu_physaddr ^ 40'h3000; // @[Parameters.scala 121:31]
  assign _T_367 = {1'b0,$signed(_T_366)}; // @[Parameters.scala 121:49]
  assign _T_369 = $signed(_T_367) & -41'sh1000; // @[Parameters.scala 121:52]
  assign _T_370 = $signed(_T_369) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_371 = mpu_physaddr ^ 40'hc000000; // @[Parameters.scala 121:31]
  assign _T_372 = {1'b0,$signed(_T_371)}; // @[Parameters.scala 121:49]
  assign _T_374 = $signed(_T_372) & -41'sh4000000; // @[Parameters.scala 121:52]
  assign _T_375 = $signed(_T_374) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_376 = mpu_physaddr ^ 40'h2000000; // @[Parameters.scala 121:31]
  assign _T_377 = {1'b0,$signed(_T_376)}; // @[Parameters.scala 121:49]
  assign _T_379 = $signed(_T_377) & -41'sh10000; // @[Parameters.scala 121:52]
  assign _T_380 = $signed(_T_379) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_382 = {1'b0,$signed(mpu_physaddr)}; // @[Parameters.scala 121:49]
  assign _T_384 = $signed(_T_382) & -41'sh1000; // @[Parameters.scala 121:52]
  assign _T_385 = $signed(_T_384) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_386 = mpu_physaddr ^ 40'h10000; // @[Parameters.scala 121:31]
  assign _T_387 = {1'b0,$signed(_T_386)}; // @[Parameters.scala 121:49]
  assign _T_389 = $signed(_T_387) & -41'sh10000; // @[Parameters.scala 121:52]
  assign _T_390 = $signed(_T_389) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_391 = mpu_physaddr ^ 40'h80000000; // @[Parameters.scala 121:31]
  assign _T_392 = {1'b0,$signed(_T_391)}; // @[Parameters.scala 121:49]
  assign _T_394 = $signed(_T_392) & -41'sh10000000; // @[Parameters.scala 121:52]
  assign _T_395 = $signed(_T_394) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_396 = mpu_physaddr ^ 40'h60000000; // @[Parameters.scala 121:31]
  assign _T_397 = {1'b0,$signed(_T_396)}; // @[Parameters.scala 121:49]
  assign _T_399 = $signed(_T_397) & -41'sh20000000; // @[Parameters.scala 121:52]
  assign _T_400 = $signed(_T_399) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_414 = _T_370 | _T_375; // @[TLB.scala 195:67]
  assign _T_415 = _T_414 | _T_380; // @[TLB.scala 195:67]
  assign _T_416 = _T_415 | _T_385; // @[TLB.scala 195:67]
  assign _T_417 = _T_416 | _T_390; // @[TLB.scala 195:67]
  assign _T_418 = _T_417 | _T_395; // @[TLB.scala 195:67]
  assign legal_address = _T_418 | _T_400; // @[TLB.scala 195:67]
  assign _T_427 = $signed(_T_392) & 41'sh80000000; // @[Parameters.scala 121:52]
  assign _T_428 = $signed(_T_427) == 41'sh0; // @[Parameters.scala 121:67]
  assign cacheable = legal_address & _T_428; // @[TLB.scala 197:19]
  assign _T_485 = mpu_physaddr ^ 40'h8000000; // @[Parameters.scala 121:31]
  assign _T_486 = {1'b0,$signed(_T_485)}; // @[Parameters.scala 121:49]
  assign _T_488 = $signed(_T_486) & 41'shc8000000; // @[Parameters.scala 121:52]
  assign _T_489 = $signed(_T_488) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_507 = $signed(_T_382) & 41'shc8010000; // @[Parameters.scala 121:52]
  assign _T_508 = $signed(_T_507) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_515 = _T_508 | _T_489; // @[TLBPermissions.scala 81:66]
  assign prot_r = legal_address & pmp_io_r; // @[TLB.scala 200:41]
  assign _T_552 = $signed(_T_392) & 41'shc0000000; // @[Parameters.scala 121:52]
  assign _T_553 = $signed(_T_552) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_554 = mpu_physaddr ^ 40'h40000000; // @[Parameters.scala 121:31]
  assign _T_555 = {1'b0,$signed(_T_554)}; // @[Parameters.scala 121:49]
  assign _T_557 = $signed(_T_555) & 41'shc0000000; // @[Parameters.scala 121:52]
  assign _T_558 = $signed(_T_557) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_560 = _T_515 | _T_553; // @[Parameters.scala 148:89]
  assign _T_561 = _T_560 | _T_558; // @[Parameters.scala 148:89]
  assign _T_568 = legal_address & _T_561; // @[TLB.scala 197:19]
  assign prot_w = _T_568 & pmp_io_w; // @[TLB.scala 201:45]
  assign _T_603 = legal_address & _T_515; // @[TLB.scala 197:19]
  assign prot_al = _T_603 | cacheable; // @[TLB.scala 202:46]
  assign _T_655 = $signed(_T_382) & 41'shca000000; // @[Parameters.scala 121:52]
  assign _T_656 = $signed(_T_655) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_667 = _T_656 | _T_553; // @[Parameters.scala 148:89]
  assign _T_668 = _T_667 | _T_558; // @[Parameters.scala 148:89]
  assign _T_675 = legal_address & _T_668; // @[TLB.scala 197:19]
  assign prot_x = _T_675 & pmp_io_x; // @[TLB.scala 204:40]
  assign _T_701 = $signed(_T_377) & 41'shca010000; // @[Parameters.scala 121:52]
  assign _T_702 = $signed(_T_701) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_706 = $signed(_T_382) & 41'shca012000; // @[Parameters.scala 121:52]
  assign _T_707 = $signed(_T_706) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_713 = _T_489 | _T_702; // @[Parameters.scala 148:89]
  assign _T_714 = _T_713 | _T_707; // @[Parameters.scala 148:89]
  assign _T_715 = _T_714 | _T_558; // @[Parameters.scala 148:89]
  assign prot_eff = legal_address & _T_715; // @[TLB.scala 197:19]
  assign _T_722 = sectored_entries_0_valid_0 | sectored_entries_0_valid_1; // @[package.scala 63:59]
  assign _T_723 = _T_722 | sectored_entries_0_valid_2; // @[package.scala 63:59]
  assign _T_724 = _T_723 | sectored_entries_0_valid_3; // @[package.scala 63:59]
  assign _T_725 = sectored_entries_0_tag ^ vpn; // @[TLB.scala 103:43]
  assign _T_727 = _T_725[26:2] == 25'h0; // @[TLB.scala 103:68]
  assign sector_hits_0 = _T_724 & _T_727; // @[TLB.scala 102:42]
  assign _T_728 = sectored_entries_1_valid_0 | sectored_entries_1_valid_1; // @[package.scala 63:59]
  assign _T_729 = _T_728 | sectored_entries_1_valid_2; // @[package.scala 63:59]
  assign _T_730 = _T_729 | sectored_entries_1_valid_3; // @[package.scala 63:59]
  assign _T_731 = sectored_entries_1_tag ^ vpn; // @[TLB.scala 103:43]
  assign _T_733 = _T_731[26:2] == 25'h0; // @[TLB.scala 103:68]
  assign sector_hits_1 = _T_730 & _T_733; // @[TLB.scala 102:42]
  assign _T_734 = sectored_entries_2_valid_0 | sectored_entries_2_valid_1; // @[package.scala 63:59]
  assign _T_735 = _T_734 | sectored_entries_2_valid_2; // @[package.scala 63:59]
  assign _T_736 = _T_735 | sectored_entries_2_valid_3; // @[package.scala 63:59]
  assign _T_737 = sectored_entries_2_tag ^ vpn; // @[TLB.scala 103:43]
  assign _T_739 = _T_737[26:2] == 25'h0; // @[TLB.scala 103:68]
  assign sector_hits_2 = _T_736 & _T_739; // @[TLB.scala 102:42]
  assign _T_740 = sectored_entries_3_valid_0 | sectored_entries_3_valid_1; // @[package.scala 63:59]
  assign _T_741 = _T_740 | sectored_entries_3_valid_2; // @[package.scala 63:59]
  assign _T_742 = _T_741 | sectored_entries_3_valid_3; // @[package.scala 63:59]
  assign _T_743 = sectored_entries_3_tag ^ vpn; // @[TLB.scala 103:43]
  assign _T_745 = _T_743[26:2] == 25'h0; // @[TLB.scala 103:68]
  assign sector_hits_3 = _T_742 & _T_745; // @[TLB.scala 102:42]
  assign _T_746 = sectored_entries_4_valid_0 | sectored_entries_4_valid_1; // @[package.scala 63:59]
  assign _T_747 = _T_746 | sectored_entries_4_valid_2; // @[package.scala 63:59]
  assign _T_748 = _T_747 | sectored_entries_4_valid_3; // @[package.scala 63:59]
  assign _T_749 = sectored_entries_4_tag ^ vpn; // @[TLB.scala 103:43]
  assign _T_751 = _T_749[26:2] == 25'h0; // @[TLB.scala 103:68]
  assign sector_hits_4 = _T_748 & _T_751; // @[TLB.scala 102:42]
  assign _T_752 = sectored_entries_5_valid_0 | sectored_entries_5_valid_1; // @[package.scala 63:59]
  assign _T_753 = _T_752 | sectored_entries_5_valid_2; // @[package.scala 63:59]
  assign _T_754 = _T_753 | sectored_entries_5_valid_3; // @[package.scala 63:59]
  assign _T_755 = sectored_entries_5_tag ^ vpn; // @[TLB.scala 103:43]
  assign _T_757 = _T_755[26:2] == 25'h0; // @[TLB.scala 103:68]
  assign sector_hits_5 = _T_754 & _T_757; // @[TLB.scala 102:42]
  assign _T_758 = sectored_entries_6_valid_0 | sectored_entries_6_valid_1; // @[package.scala 63:59]
  assign _T_759 = _T_758 | sectored_entries_6_valid_2; // @[package.scala 63:59]
  assign _T_760 = _T_759 | sectored_entries_6_valid_3; // @[package.scala 63:59]
  assign _T_761 = sectored_entries_6_tag ^ vpn; // @[TLB.scala 103:43]
  assign _T_763 = _T_761[26:2] == 25'h0; // @[TLB.scala 103:68]
  assign sector_hits_6 = _T_760 & _T_763; // @[TLB.scala 102:42]
  assign _T_764 = sectored_entries_7_valid_0 | sectored_entries_7_valid_1; // @[package.scala 63:59]
  assign _T_765 = _T_764 | sectored_entries_7_valid_2; // @[package.scala 63:59]
  assign _T_766 = _T_765 | sectored_entries_7_valid_3; // @[package.scala 63:59]
  assign _T_767 = sectored_entries_7_tag ^ vpn; // @[TLB.scala 103:43]
  assign _T_769 = _T_767[26:2] == 25'h0; // @[TLB.scala 103:68]
  assign sector_hits_7 = _T_766 & _T_769; // @[TLB.scala 102:42]
  assign _T_774 = superpage_entries_0_tag[26:18] == vpn[26:18]; // @[TLB.scala 110:79]
  assign _T_776 = superpage_entries_0_valid_0 & _T_774; // @[TLB.scala 110:31]
  assign _T_777 = superpage_entries_0_level < 2'h1; // @[TLB.scala 109:30]
  assign _T_781 = superpage_entries_0_tag[17:9] == vpn[17:9]; // @[TLB.scala 110:79]
  assign _T_782 = _T_777 | _T_781; // @[TLB.scala 110:42]
  assign superpage_hits_0 = _T_776 & _T_782; // @[TLB.scala 110:31]
  assign _T_794 = superpage_entries_1_tag[26:18] == vpn[26:18]; // @[TLB.scala 110:79]
  assign _T_796 = superpage_entries_1_valid_0 & _T_794; // @[TLB.scala 110:31]
  assign _T_797 = superpage_entries_1_level < 2'h1; // @[TLB.scala 109:30]
  assign _T_801 = superpage_entries_1_tag[17:9] == vpn[17:9]; // @[TLB.scala 110:79]
  assign _T_802 = _T_797 | _T_801; // @[TLB.scala 110:42]
  assign superpage_hits_1 = _T_796 & _T_802; // @[TLB.scala 110:31]
  assign _T_814 = superpage_entries_2_tag[26:18] == vpn[26:18]; // @[TLB.scala 110:79]
  assign _T_816 = superpage_entries_2_valid_0 & _T_814; // @[TLB.scala 110:31]
  assign _T_817 = superpage_entries_2_level < 2'h1; // @[TLB.scala 109:30]
  assign _T_821 = superpage_entries_2_tag[17:9] == vpn[17:9]; // @[TLB.scala 110:79]
  assign _T_822 = _T_817 | _T_821; // @[TLB.scala 110:42]
  assign superpage_hits_2 = _T_816 & _T_822; // @[TLB.scala 110:31]
  assign _T_834 = superpage_entries_3_tag[26:18] == vpn[26:18]; // @[TLB.scala 110:79]
  assign _T_836 = superpage_entries_3_valid_0 & _T_834; // @[TLB.scala 110:31]
  assign _T_837 = superpage_entries_3_level < 2'h1; // @[TLB.scala 109:30]
  assign _T_841 = superpage_entries_3_tag[17:9] == vpn[17:9]; // @[TLB.scala 110:79]
  assign _T_842 = _T_837 | _T_841; // @[TLB.scala 110:42]
  assign superpage_hits_3 = _T_836 & _T_842; // @[TLB.scala 110:31]
  assign _GEN_1 = 2'h1 == vpn[1:0] ? sectored_entries_0_valid_1 : sectored_entries_0_valid_0; // @[TLB.scala 115:20]
  assign _GEN_2 = 2'h2 == vpn[1:0] ? sectored_entries_0_valid_2 : _GEN_1; // @[TLB.scala 115:20]
  assign _GEN_3 = 2'h3 == vpn[1:0] ? sectored_entries_0_valid_3 : _GEN_2; // @[TLB.scala 115:20]
  assign _T_854 = _GEN_3 & _T_727; // @[TLB.scala 115:20]
  assign hitsVec_0 = vm_enabled & _T_854; // @[TLB.scala 209:44]
  assign _GEN_5 = 2'h1 == vpn[1:0] ? sectored_entries_1_valid_1 : sectored_entries_1_valid_0; // @[TLB.scala 115:20]
  assign _GEN_6 = 2'h2 == vpn[1:0] ? sectored_entries_1_valid_2 : _GEN_5; // @[TLB.scala 115:20]
  assign _GEN_7 = 2'h3 == vpn[1:0] ? sectored_entries_1_valid_3 : _GEN_6; // @[TLB.scala 115:20]
  assign _T_859 = _GEN_7 & _T_733; // @[TLB.scala 115:20]
  assign hitsVec_1 = vm_enabled & _T_859; // @[TLB.scala 209:44]
  assign _GEN_9 = 2'h1 == vpn[1:0] ? sectored_entries_2_valid_1 : sectored_entries_2_valid_0; // @[TLB.scala 115:20]
  assign _GEN_10 = 2'h2 == vpn[1:0] ? sectored_entries_2_valid_2 : _GEN_9; // @[TLB.scala 115:20]
  assign _GEN_11 = 2'h3 == vpn[1:0] ? sectored_entries_2_valid_3 : _GEN_10; // @[TLB.scala 115:20]
  assign _T_864 = _GEN_11 & _T_739; // @[TLB.scala 115:20]
  assign hitsVec_2 = vm_enabled & _T_864; // @[TLB.scala 209:44]
  assign _GEN_13 = 2'h1 == vpn[1:0] ? sectored_entries_3_valid_1 : sectored_entries_3_valid_0; // @[TLB.scala 115:20]
  assign _GEN_14 = 2'h2 == vpn[1:0] ? sectored_entries_3_valid_2 : _GEN_13; // @[TLB.scala 115:20]
  assign _GEN_15 = 2'h3 == vpn[1:0] ? sectored_entries_3_valid_3 : _GEN_14; // @[TLB.scala 115:20]
  assign _T_869 = _GEN_15 & _T_745; // @[TLB.scala 115:20]
  assign hitsVec_3 = vm_enabled & _T_869; // @[TLB.scala 209:44]
  assign _GEN_17 = 2'h1 == vpn[1:0] ? sectored_entries_4_valid_1 : sectored_entries_4_valid_0; // @[TLB.scala 115:20]
  assign _GEN_18 = 2'h2 == vpn[1:0] ? sectored_entries_4_valid_2 : _GEN_17; // @[TLB.scala 115:20]
  assign _GEN_19 = 2'h3 == vpn[1:0] ? sectored_entries_4_valid_3 : _GEN_18; // @[TLB.scala 115:20]
  assign _T_874 = _GEN_19 & _T_751; // @[TLB.scala 115:20]
  assign hitsVec_4 = vm_enabled & _T_874; // @[TLB.scala 209:44]
  assign _GEN_21 = 2'h1 == vpn[1:0] ? sectored_entries_5_valid_1 : sectored_entries_5_valid_0; // @[TLB.scala 115:20]
  assign _GEN_22 = 2'h2 == vpn[1:0] ? sectored_entries_5_valid_2 : _GEN_21; // @[TLB.scala 115:20]
  assign _GEN_23 = 2'h3 == vpn[1:0] ? sectored_entries_5_valid_3 : _GEN_22; // @[TLB.scala 115:20]
  assign _T_879 = _GEN_23 & _T_757; // @[TLB.scala 115:20]
  assign hitsVec_5 = vm_enabled & _T_879; // @[TLB.scala 209:44]
  assign _GEN_25 = 2'h1 == vpn[1:0] ? sectored_entries_6_valid_1 : sectored_entries_6_valid_0; // @[TLB.scala 115:20]
  assign _GEN_26 = 2'h2 == vpn[1:0] ? sectored_entries_6_valid_2 : _GEN_25; // @[TLB.scala 115:20]
  assign _GEN_27 = 2'h3 == vpn[1:0] ? sectored_entries_6_valid_3 : _GEN_26; // @[TLB.scala 115:20]
  assign _T_884 = _GEN_27 & _T_763; // @[TLB.scala 115:20]
  assign hitsVec_6 = vm_enabled & _T_884; // @[TLB.scala 209:44]
  assign _GEN_29 = 2'h1 == vpn[1:0] ? sectored_entries_7_valid_1 : sectored_entries_7_valid_0; // @[TLB.scala 115:20]
  assign _GEN_30 = 2'h2 == vpn[1:0] ? sectored_entries_7_valid_2 : _GEN_29; // @[TLB.scala 115:20]
  assign _GEN_31 = 2'h3 == vpn[1:0] ? sectored_entries_7_valid_3 : _GEN_30; // @[TLB.scala 115:20]
  assign _T_889 = _GEN_31 & _T_769; // @[TLB.scala 115:20]
  assign hitsVec_7 = vm_enabled & _T_889; // @[TLB.scala 209:44]
  assign hitsVec_8 = vm_enabled & superpage_hits_0; // @[TLB.scala 209:44]
  assign hitsVec_9 = vm_enabled & superpage_hits_1; // @[TLB.scala 209:44]
  assign hitsVec_10 = vm_enabled & superpage_hits_2; // @[TLB.scala 209:44]
  assign hitsVec_11 = vm_enabled & superpage_hits_3; // @[TLB.scala 209:44]
  assign _T_978 = special_entry_tag[26:18] == vpn[26:18]; // @[TLB.scala 110:79]
  assign _T_980 = special_entry_valid_0 & _T_978; // @[TLB.scala 110:31]
  assign _T_985 = special_entry_tag[17:9] == vpn[17:9]; // @[TLB.scala 110:79]
  assign _T_986 = _T_348 | _T_985; // @[TLB.scala 110:42]
  assign _T_987 = _T_980 & _T_986; // @[TLB.scala 110:31]
  assign _T_992 = special_entry_tag[8:0] == vpn[8:0]; // @[TLB.scala 110:79]
  assign _T_993 = _T_354 | _T_992; // @[TLB.scala 110:42]
  assign _T_994 = _T_987 & _T_993; // @[TLB.scala 110:31]
  assign hitsVec_12 = vm_enabled & _T_994; // @[TLB.scala 209:44]
  assign _T_999 = {hitsVec_5,hitsVec_4,hitsVec_3,hitsVec_2,hitsVec_1,hitsVec_0}; // @[Cat.scala 30:58]
  assign real_hits = {hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,_T_999}; // @[Cat.scala 30:58]
  assign hits = {~vm_enabled,hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,_T_999}; // @[Cat.scala 30:58]
  assign _GEN_33 = 2'h1 == vpn[1:0] ? sectored_entries_0_data_1 : sectored_entries_0_data_0;
  assign _GEN_34 = 2'h2 == vpn[1:0] ? sectored_entries_0_data_2 : _GEN_33;
  assign _GEN_35 = 2'h3 == vpn[1:0] ? sectored_entries_0_data_3 : _GEN_34;
  assign _GEN_37 = 2'h1 == vpn[1:0] ? sectored_entries_1_data_1 : sectored_entries_1_data_0;
  assign _GEN_38 = 2'h2 == vpn[1:0] ? sectored_entries_1_data_2 : _GEN_37;
  assign _GEN_39 = 2'h3 == vpn[1:0] ? sectored_entries_1_data_3 : _GEN_38;
  assign _GEN_41 = 2'h1 == vpn[1:0] ? sectored_entries_2_data_1 : sectored_entries_2_data_0;
  assign _GEN_42 = 2'h2 == vpn[1:0] ? sectored_entries_2_data_2 : _GEN_41;
  assign _GEN_43 = 2'h3 == vpn[1:0] ? sectored_entries_2_data_3 : _GEN_42;
  assign _GEN_45 = 2'h1 == vpn[1:0] ? sectored_entries_3_data_1 : sectored_entries_3_data_0;
  assign _GEN_46 = 2'h2 == vpn[1:0] ? sectored_entries_3_data_2 : _GEN_45;
  assign _GEN_47 = 2'h3 == vpn[1:0] ? sectored_entries_3_data_3 : _GEN_46;
  assign _GEN_49 = 2'h1 == vpn[1:0] ? sectored_entries_4_data_1 : sectored_entries_4_data_0;
  assign _GEN_50 = 2'h2 == vpn[1:0] ? sectored_entries_4_data_2 : _GEN_49;
  assign _GEN_51 = 2'h3 == vpn[1:0] ? sectored_entries_4_data_3 : _GEN_50;
  assign _GEN_53 = 2'h1 == vpn[1:0] ? sectored_entries_5_data_1 : sectored_entries_5_data_0;
  assign _GEN_54 = 2'h2 == vpn[1:0] ? sectored_entries_5_data_2 : _GEN_53;
  assign _GEN_55 = 2'h3 == vpn[1:0] ? sectored_entries_5_data_3 : _GEN_54;
  assign _GEN_57 = 2'h1 == vpn[1:0] ? sectored_entries_6_data_1 : sectored_entries_6_data_0;
  assign _GEN_58 = 2'h2 == vpn[1:0] ? sectored_entries_6_data_2 : _GEN_57;
  assign _GEN_59 = 2'h3 == vpn[1:0] ? sectored_entries_6_data_3 : _GEN_58;
  assign _GEN_61 = 2'h1 == vpn[1:0] ? sectored_entries_7_data_1 : sectored_entries_7_data_0;
  assign _GEN_62 = 2'h2 == vpn[1:0] ? sectored_entries_7_data_2 : _GEN_61;
  assign _GEN_63 = 2'h3 == vpn[1:0] ? sectored_entries_7_data_3 : _GEN_62;
  assign _T_1199 = _T_777 ? vpn : 27'h0; // @[TLB.scala 124:30]
  assign _GEN_956 = {{7'd0}, superpage_entries_0_data_0[33:14]}; // @[TLB.scala 124:49]
  assign _T_1200 = _T_1199 | _GEN_956; // @[TLB.scala 124:49]
  assign _T_1206 = vpn | _GEN_956; // @[TLB.scala 124:49]
  assign _T_1208 = {superpage_entries_0_data_0[33:32],_T_1200[17:9],_T_1206[8:0]}; // @[Cat.scala 30:58]
  assign _T_1232 = _T_797 ? vpn : 27'h0; // @[TLB.scala 124:30]
  assign _GEN_958 = {{7'd0}, superpage_entries_1_data_0[33:14]}; // @[TLB.scala 124:49]
  assign _T_1233 = _T_1232 | _GEN_958; // @[TLB.scala 124:49]
  assign _T_1239 = vpn | _GEN_958; // @[TLB.scala 124:49]
  assign _T_1241 = {superpage_entries_1_data_0[33:32],_T_1233[17:9],_T_1239[8:0]}; // @[Cat.scala 30:58]
  assign _T_1265 = _T_817 ? vpn : 27'h0; // @[TLB.scala 124:30]
  assign _GEN_960 = {{7'd0}, superpage_entries_2_data_0[33:14]}; // @[TLB.scala 124:49]
  assign _T_1266 = _T_1265 | _GEN_960; // @[TLB.scala 124:49]
  assign _T_1272 = vpn | _GEN_960; // @[TLB.scala 124:49]
  assign _T_1274 = {superpage_entries_2_data_0[33:32],_T_1266[17:9],_T_1272[8:0]}; // @[Cat.scala 30:58]
  assign _T_1298 = _T_837 ? vpn : 27'h0; // @[TLB.scala 124:30]
  assign _GEN_962 = {{7'd0}, superpage_entries_3_data_0[33:14]}; // @[TLB.scala 124:49]
  assign _T_1299 = _T_1298 | _GEN_962; // @[TLB.scala 124:49]
  assign _T_1305 = vpn | _GEN_962; // @[TLB.scala 124:49]
  assign _T_1307 = {superpage_entries_3_data_0[33:32],_T_1299[17:9],_T_1305[8:0]}; // @[Cat.scala 30:58]
  assign _T_1343 = hitsVec_0 ? _GEN_35[33:14] : 20'h0; // @[Mux.scala 19:72]
  assign _T_1344 = hitsVec_1 ? _GEN_39[33:14] : 20'h0; // @[Mux.scala 19:72]
  assign _T_1345 = hitsVec_2 ? _GEN_43[33:14] : 20'h0; // @[Mux.scala 19:72]
  assign _T_1346 = hitsVec_3 ? _GEN_47[33:14] : 20'h0; // @[Mux.scala 19:72]
  assign _T_1347 = hitsVec_4 ? _GEN_51[33:14] : 20'h0; // @[Mux.scala 19:72]
  assign _T_1348 = hitsVec_5 ? _GEN_55[33:14] : 20'h0; // @[Mux.scala 19:72]
  assign _T_1349 = hitsVec_6 ? _GEN_59[33:14] : 20'h0; // @[Mux.scala 19:72]
  assign _T_1350 = hitsVec_7 ? _GEN_63[33:14] : 20'h0; // @[Mux.scala 19:72]
  assign _T_1351 = hitsVec_8 ? _T_1208 : 20'h0; // @[Mux.scala 19:72]
  assign _T_1352 = hitsVec_9 ? _T_1241 : 20'h0; // @[Mux.scala 19:72]
  assign _T_1353 = hitsVec_10 ? _T_1274 : 20'h0; // @[Mux.scala 19:72]
  assign _T_1354 = hitsVec_11 ? _T_1307 : 20'h0; // @[Mux.scala 19:72]
  assign _T_1355 = hitsVec_12 ? _T_359 : 20'h0; // @[Mux.scala 19:72]
  assign _T_1356 = vm_enabled ? 20'h0 : vpn[19:0]; // @[Mux.scala 19:72]
  assign _T_1357 = _T_1343 | _T_1344; // @[Mux.scala 19:72]
  assign _T_1358 = _T_1357 | _T_1345; // @[Mux.scala 19:72]
  assign _T_1359 = _T_1358 | _T_1346; // @[Mux.scala 19:72]
  assign _T_1360 = _T_1359 | _T_1347; // @[Mux.scala 19:72]
  assign _T_1361 = _T_1360 | _T_1348; // @[Mux.scala 19:72]
  assign _T_1362 = _T_1361 | _T_1349; // @[Mux.scala 19:72]
  assign _T_1363 = _T_1362 | _T_1350; // @[Mux.scala 19:72]
  assign _T_1364 = _T_1363 | _T_1351; // @[Mux.scala 19:72]
  assign _T_1365 = _T_1364 | _T_1352; // @[Mux.scala 19:72]
  assign _T_1366 = _T_1365 | _T_1353; // @[Mux.scala 19:72]
  assign _T_1367 = _T_1366 | _T_1354; // @[Mux.scala 19:72]
  assign _T_1368 = _T_1367 | _T_1355; // @[Mux.scala 19:72]
  assign ppn = _T_1368 | _T_1356; // @[Mux.scala 19:72]
  assign _T_1385 = io_ptw_resp_valid & ~invalidate_refill; // @[TLB.scala 224:17]
  assign _GEN_966 = {{27'd0}, vpoffset_cfg_value}; // @[TLB.scala 227:31]
  assign _T_1387 = io_ptw_resp_bits_pte_ppn + _GEN_966; // @[TLB.scala 227:31]
  assign _T_1391 = io_ptw_resp_bits_pte_x & ~io_ptw_resp_bits_pte_w; // @[PTW.scala 77:44]
  assign _T_1392 = io_ptw_resp_bits_pte_r | _T_1391; // @[PTW.scala 77:38]
  assign _T_1393 = io_ptw_resp_bits_pte_v & _T_1392; // @[PTW.scala 77:32]
  assign _T_1394 = _T_1393 & io_ptw_resp_bits_pte_a; // @[PTW.scala 77:52]
  assign _T_1395 = _T_1394 & io_ptw_resp_bits_pte_r; // @[PTW.scala 81:35]
  assign _T_1401 = _T_1394 & io_ptw_resp_bits_pte_w; // @[PTW.scala 82:35]
  assign _T_1402 = _T_1401 & io_ptw_resp_bits_pte_d; // @[PTW.scala 82:40]
  assign _T_1403 = vpoffset_cfg_value == 27'h0; // @[TLB.scala 231:55]
  assign _T_1404 = io_ptw_resp_bits_pte_u | _T_1403; // @[TLB.scala 231:32]
  assign _T_1405 = io_ptw_resp_bits_level != 2'h2; // @[TLB.scala 231:90]
  assign _T_1406 = _T_1404 | _T_1405; // @[TLB.scala 231:64]
  assign _T_1412 = _T_1394 & io_ptw_resp_bits_pte_x; // @[PTW.scala 83:35]
  assign _GEN_967 = {{27'd0}, requestedVPN}; // @[TLB.scala 231:133]
  assign _T_1413 = _T_1387 == _GEN_967; // @[TLB.scala 231:133]
  assign _T_1420 = _T_1413 & _T_1412; // @[TLB.scala 231:120]
  assign _T_1421 = _T_1406 ? _T_1412 : _T_1420; // @[TLB.scala 231:25]
  assign _T_1430 = {prot_x,prot_r,prot_al,prot_al,prot_eff,cacheable,1'h0}; // @[TLB.scala 138:26]
  assign _T_1438 = {refill_ppn,io_ptw_resp_bits_pte_u,io_ptw_resp_bits_pte_g,io_ptw_resp_bits_ae,_T_1402,_T_1421,_T_1395,prot_w,_T_1430}; // @[TLB.scala 138:26]
  assign _T_1439 = io_ptw_resp_bits_level < 2'h2; // @[TLB.scala 253:40]
  assign _T_1440 = r_superpage_repl_addr == 2'h0; // @[TLB.scala 254:82]
  assign _GEN_67 = _T_1440 | superpage_entries_0_valid_0; // @[TLB.scala 254:89]
  assign _T_1456 = r_superpage_repl_addr == 2'h1; // @[TLB.scala 254:82]
  assign _GEN_71 = _T_1456 | superpage_entries_1_valid_0; // @[TLB.scala 254:89]
  assign _T_1472 = r_superpage_repl_addr == 2'h2; // @[TLB.scala 254:82]
  assign _GEN_75 = _T_1472 | superpage_entries_2_valid_0; // @[TLB.scala 254:89]
  assign _T_1488 = r_superpage_repl_addr == 2'h3; // @[TLB.scala 254:82]
  assign _GEN_79 = _T_1488 | superpage_entries_3_valid_0; // @[TLB.scala 254:89]
  assign _T_1504 = r_sectored_hit ? r_sectored_hit_addr : r_sectored_repl_addr; // @[TLB.scala 258:22]
  assign _T_1505 = _T_1504 == 3'h0; // @[TLB.scala 259:65]
  assign _GEN_81 = r_sectored_hit ? sectored_entries_0_valid_0 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_82 = r_sectored_hit ? sectored_entries_0_valid_1 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_83 = r_sectored_hit ? sectored_entries_0_valid_2 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_84 = r_sectored_hit ? sectored_entries_0_valid_3 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_968 = 2'h0 == r_refill_tag[1:0]; // @[TLB.scala 137:18]
  assign _GEN_85 = _GEN_968 | _GEN_81; // @[TLB.scala 137:18]
  assign _GEN_969 = 2'h1 == r_refill_tag[1:0]; // @[TLB.scala 137:18]
  assign _GEN_86 = _GEN_969 | _GEN_82; // @[TLB.scala 137:18]
  assign _GEN_970 = 2'h2 == r_refill_tag[1:0]; // @[TLB.scala 137:18]
  assign _GEN_87 = _GEN_970 | _GEN_83; // @[TLB.scala 137:18]
  assign _GEN_971 = 2'h3 == r_refill_tag[1:0]; // @[TLB.scala 137:18]
  assign _GEN_88 = _GEN_971 | _GEN_84; // @[TLB.scala 137:18]
  assign _GEN_93 = _T_1505 ? _GEN_85 : sectored_entries_0_valid_0; // @[TLB.scala 259:72]
  assign _GEN_94 = _T_1505 ? _GEN_86 : sectored_entries_0_valid_1; // @[TLB.scala 259:72]
  assign _GEN_95 = _T_1505 ? _GEN_87 : sectored_entries_0_valid_2; // @[TLB.scala 259:72]
  assign _GEN_96 = _T_1505 ? _GEN_88 : sectored_entries_0_valid_3; // @[TLB.scala 259:72]
  assign _T_1522 = _T_1504 == 3'h1; // @[TLB.scala 259:65]
  assign _GEN_103 = r_sectored_hit ? sectored_entries_1_valid_0 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_104 = r_sectored_hit ? sectored_entries_1_valid_1 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_105 = r_sectored_hit ? sectored_entries_1_valid_2 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_106 = r_sectored_hit ? sectored_entries_1_valid_3 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_107 = _GEN_968 | _GEN_103; // @[TLB.scala 137:18]
  assign _GEN_108 = _GEN_969 | _GEN_104; // @[TLB.scala 137:18]
  assign _GEN_109 = _GEN_970 | _GEN_105; // @[TLB.scala 137:18]
  assign _GEN_110 = _GEN_971 | _GEN_106; // @[TLB.scala 137:18]
  assign _GEN_115 = _T_1522 ? _GEN_107 : sectored_entries_1_valid_0; // @[TLB.scala 259:72]
  assign _GEN_116 = _T_1522 ? _GEN_108 : sectored_entries_1_valid_1; // @[TLB.scala 259:72]
  assign _GEN_117 = _T_1522 ? _GEN_109 : sectored_entries_1_valid_2; // @[TLB.scala 259:72]
  assign _GEN_118 = _T_1522 ? _GEN_110 : sectored_entries_1_valid_3; // @[TLB.scala 259:72]
  assign _T_1539 = _T_1504 == 3'h2; // @[TLB.scala 259:65]
  assign _GEN_125 = r_sectored_hit ? sectored_entries_2_valid_0 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_126 = r_sectored_hit ? sectored_entries_2_valid_1 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_127 = r_sectored_hit ? sectored_entries_2_valid_2 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_128 = r_sectored_hit ? sectored_entries_2_valid_3 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_129 = _GEN_968 | _GEN_125; // @[TLB.scala 137:18]
  assign _GEN_130 = _GEN_969 | _GEN_126; // @[TLB.scala 137:18]
  assign _GEN_131 = _GEN_970 | _GEN_127; // @[TLB.scala 137:18]
  assign _GEN_132 = _GEN_971 | _GEN_128; // @[TLB.scala 137:18]
  assign _GEN_137 = _T_1539 ? _GEN_129 : sectored_entries_2_valid_0; // @[TLB.scala 259:72]
  assign _GEN_138 = _T_1539 ? _GEN_130 : sectored_entries_2_valid_1; // @[TLB.scala 259:72]
  assign _GEN_139 = _T_1539 ? _GEN_131 : sectored_entries_2_valid_2; // @[TLB.scala 259:72]
  assign _GEN_140 = _T_1539 ? _GEN_132 : sectored_entries_2_valid_3; // @[TLB.scala 259:72]
  assign _T_1556 = _T_1504 == 3'h3; // @[TLB.scala 259:65]
  assign _GEN_147 = r_sectored_hit ? sectored_entries_3_valid_0 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_148 = r_sectored_hit ? sectored_entries_3_valid_1 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_149 = r_sectored_hit ? sectored_entries_3_valid_2 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_150 = r_sectored_hit ? sectored_entries_3_valid_3 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_151 = _GEN_968 | _GEN_147; // @[TLB.scala 137:18]
  assign _GEN_152 = _GEN_969 | _GEN_148; // @[TLB.scala 137:18]
  assign _GEN_153 = _GEN_970 | _GEN_149; // @[TLB.scala 137:18]
  assign _GEN_154 = _GEN_971 | _GEN_150; // @[TLB.scala 137:18]
  assign _GEN_159 = _T_1556 ? _GEN_151 : sectored_entries_3_valid_0; // @[TLB.scala 259:72]
  assign _GEN_160 = _T_1556 ? _GEN_152 : sectored_entries_3_valid_1; // @[TLB.scala 259:72]
  assign _GEN_161 = _T_1556 ? _GEN_153 : sectored_entries_3_valid_2; // @[TLB.scala 259:72]
  assign _GEN_162 = _T_1556 ? _GEN_154 : sectored_entries_3_valid_3; // @[TLB.scala 259:72]
  assign _T_1573 = _T_1504 == 3'h4; // @[TLB.scala 259:65]
  assign _GEN_169 = r_sectored_hit ? sectored_entries_4_valid_0 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_170 = r_sectored_hit ? sectored_entries_4_valid_1 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_171 = r_sectored_hit ? sectored_entries_4_valid_2 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_172 = r_sectored_hit ? sectored_entries_4_valid_3 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_173 = _GEN_968 | _GEN_169; // @[TLB.scala 137:18]
  assign _GEN_174 = _GEN_969 | _GEN_170; // @[TLB.scala 137:18]
  assign _GEN_175 = _GEN_970 | _GEN_171; // @[TLB.scala 137:18]
  assign _GEN_176 = _GEN_971 | _GEN_172; // @[TLB.scala 137:18]
  assign _GEN_181 = _T_1573 ? _GEN_173 : sectored_entries_4_valid_0; // @[TLB.scala 259:72]
  assign _GEN_182 = _T_1573 ? _GEN_174 : sectored_entries_4_valid_1; // @[TLB.scala 259:72]
  assign _GEN_183 = _T_1573 ? _GEN_175 : sectored_entries_4_valid_2; // @[TLB.scala 259:72]
  assign _GEN_184 = _T_1573 ? _GEN_176 : sectored_entries_4_valid_3; // @[TLB.scala 259:72]
  assign _T_1590 = _T_1504 == 3'h5; // @[TLB.scala 259:65]
  assign _GEN_191 = r_sectored_hit ? sectored_entries_5_valid_0 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_192 = r_sectored_hit ? sectored_entries_5_valid_1 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_193 = r_sectored_hit ? sectored_entries_5_valid_2 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_194 = r_sectored_hit ? sectored_entries_5_valid_3 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_195 = _GEN_968 | _GEN_191; // @[TLB.scala 137:18]
  assign _GEN_196 = _GEN_969 | _GEN_192; // @[TLB.scala 137:18]
  assign _GEN_197 = _GEN_970 | _GEN_193; // @[TLB.scala 137:18]
  assign _GEN_198 = _GEN_971 | _GEN_194; // @[TLB.scala 137:18]
  assign _GEN_203 = _T_1590 ? _GEN_195 : sectored_entries_5_valid_0; // @[TLB.scala 259:72]
  assign _GEN_204 = _T_1590 ? _GEN_196 : sectored_entries_5_valid_1; // @[TLB.scala 259:72]
  assign _GEN_205 = _T_1590 ? _GEN_197 : sectored_entries_5_valid_2; // @[TLB.scala 259:72]
  assign _GEN_206 = _T_1590 ? _GEN_198 : sectored_entries_5_valid_3; // @[TLB.scala 259:72]
  assign _T_1607 = _T_1504 == 3'h6; // @[TLB.scala 259:65]
  assign _GEN_213 = r_sectored_hit ? sectored_entries_6_valid_0 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_214 = r_sectored_hit ? sectored_entries_6_valid_1 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_215 = r_sectored_hit ? sectored_entries_6_valid_2 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_216 = r_sectored_hit ? sectored_entries_6_valid_3 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_217 = _GEN_968 | _GEN_213; // @[TLB.scala 137:18]
  assign _GEN_218 = _GEN_969 | _GEN_214; // @[TLB.scala 137:18]
  assign _GEN_219 = _GEN_970 | _GEN_215; // @[TLB.scala 137:18]
  assign _GEN_220 = _GEN_971 | _GEN_216; // @[TLB.scala 137:18]
  assign _GEN_225 = _T_1607 ? _GEN_217 : sectored_entries_6_valid_0; // @[TLB.scala 259:72]
  assign _GEN_226 = _T_1607 ? _GEN_218 : sectored_entries_6_valid_1; // @[TLB.scala 259:72]
  assign _GEN_227 = _T_1607 ? _GEN_219 : sectored_entries_6_valid_2; // @[TLB.scala 259:72]
  assign _GEN_228 = _T_1607 ? _GEN_220 : sectored_entries_6_valid_3; // @[TLB.scala 259:72]
  assign _T_1624 = _T_1504 == 3'h7; // @[TLB.scala 259:65]
  assign _GEN_235 = r_sectored_hit ? sectored_entries_7_valid_0 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_236 = r_sectored_hit ? sectored_entries_7_valid_1 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_237 = r_sectored_hit ? sectored_entries_7_valid_2 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_238 = r_sectored_hit ? sectored_entries_7_valid_3 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_239 = _GEN_968 | _GEN_235; // @[TLB.scala 137:18]
  assign _GEN_240 = _GEN_969 | _GEN_236; // @[TLB.scala 137:18]
  assign _GEN_241 = _GEN_970 | _GEN_237; // @[TLB.scala 137:18]
  assign _GEN_242 = _GEN_971 | _GEN_238; // @[TLB.scala 137:18]
  assign _GEN_247 = _T_1624 ? _GEN_239 : sectored_entries_7_valid_0; // @[TLB.scala 259:72]
  assign _GEN_248 = _T_1624 ? _GEN_240 : sectored_entries_7_valid_1; // @[TLB.scala 259:72]
  assign _GEN_249 = _T_1624 ? _GEN_241 : sectored_entries_7_valid_2; // @[TLB.scala 259:72]
  assign _GEN_250 = _T_1624 ? _GEN_242 : sectored_entries_7_valid_3; // @[TLB.scala 259:72]
  assign _GEN_259 = _T_1439 ? _GEN_67 : superpage_entries_0_valid_0; // @[TLB.scala 253:54]
  assign _GEN_263 = _T_1439 ? _GEN_71 : superpage_entries_1_valid_0; // @[TLB.scala 253:54]
  assign _GEN_267 = _T_1439 ? _GEN_75 : superpage_entries_2_valid_0; // @[TLB.scala 253:54]
  assign _GEN_271 = _T_1439 ? _GEN_79 : superpage_entries_3_valid_0; // @[TLB.scala 253:54]
  assign _GEN_273 = _T_1439 ? sectored_entries_0_valid_0 : _GEN_93; // @[TLB.scala 253:54]
  assign _GEN_274 = _T_1439 ? sectored_entries_0_valid_1 : _GEN_94; // @[TLB.scala 253:54]
  assign _GEN_275 = _T_1439 ? sectored_entries_0_valid_2 : _GEN_95; // @[TLB.scala 253:54]
  assign _GEN_276 = _T_1439 ? sectored_entries_0_valid_3 : _GEN_96; // @[TLB.scala 253:54]
  assign _GEN_283 = _T_1439 ? sectored_entries_1_valid_0 : _GEN_115; // @[TLB.scala 253:54]
  assign _GEN_284 = _T_1439 ? sectored_entries_1_valid_1 : _GEN_116; // @[TLB.scala 253:54]
  assign _GEN_285 = _T_1439 ? sectored_entries_1_valid_2 : _GEN_117; // @[TLB.scala 253:54]
  assign _GEN_286 = _T_1439 ? sectored_entries_1_valid_3 : _GEN_118; // @[TLB.scala 253:54]
  assign _GEN_293 = _T_1439 ? sectored_entries_2_valid_0 : _GEN_137; // @[TLB.scala 253:54]
  assign _GEN_294 = _T_1439 ? sectored_entries_2_valid_1 : _GEN_138; // @[TLB.scala 253:54]
  assign _GEN_295 = _T_1439 ? sectored_entries_2_valid_2 : _GEN_139; // @[TLB.scala 253:54]
  assign _GEN_296 = _T_1439 ? sectored_entries_2_valid_3 : _GEN_140; // @[TLB.scala 253:54]
  assign _GEN_303 = _T_1439 ? sectored_entries_3_valid_0 : _GEN_159; // @[TLB.scala 253:54]
  assign _GEN_304 = _T_1439 ? sectored_entries_3_valid_1 : _GEN_160; // @[TLB.scala 253:54]
  assign _GEN_305 = _T_1439 ? sectored_entries_3_valid_2 : _GEN_161; // @[TLB.scala 253:54]
  assign _GEN_306 = _T_1439 ? sectored_entries_3_valid_3 : _GEN_162; // @[TLB.scala 253:54]
  assign _GEN_313 = _T_1439 ? sectored_entries_4_valid_0 : _GEN_181; // @[TLB.scala 253:54]
  assign _GEN_314 = _T_1439 ? sectored_entries_4_valid_1 : _GEN_182; // @[TLB.scala 253:54]
  assign _GEN_315 = _T_1439 ? sectored_entries_4_valid_2 : _GEN_183; // @[TLB.scala 253:54]
  assign _GEN_316 = _T_1439 ? sectored_entries_4_valid_3 : _GEN_184; // @[TLB.scala 253:54]
  assign _GEN_323 = _T_1439 ? sectored_entries_5_valid_0 : _GEN_203; // @[TLB.scala 253:54]
  assign _GEN_324 = _T_1439 ? sectored_entries_5_valid_1 : _GEN_204; // @[TLB.scala 253:54]
  assign _GEN_325 = _T_1439 ? sectored_entries_5_valid_2 : _GEN_205; // @[TLB.scala 253:54]
  assign _GEN_326 = _T_1439 ? sectored_entries_5_valid_3 : _GEN_206; // @[TLB.scala 253:54]
  assign _GEN_333 = _T_1439 ? sectored_entries_6_valid_0 : _GEN_225; // @[TLB.scala 253:54]
  assign _GEN_334 = _T_1439 ? sectored_entries_6_valid_1 : _GEN_226; // @[TLB.scala 253:54]
  assign _GEN_335 = _T_1439 ? sectored_entries_6_valid_2 : _GEN_227; // @[TLB.scala 253:54]
  assign _GEN_336 = _T_1439 ? sectored_entries_6_valid_3 : _GEN_228; // @[TLB.scala 253:54]
  assign _GEN_343 = _T_1439 ? sectored_entries_7_valid_0 : _GEN_247; // @[TLB.scala 253:54]
  assign _GEN_344 = _T_1439 ? sectored_entries_7_valid_1 : _GEN_248; // @[TLB.scala 253:54]
  assign _GEN_345 = _T_1439 ? sectored_entries_7_valid_2 : _GEN_249; // @[TLB.scala 253:54]
  assign _GEN_346 = _T_1439 ? sectored_entries_7_valid_3 : _GEN_250; // @[TLB.scala 253:54]
  assign _GEN_355 = ~io_ptw_resp_bits_homogeneous | special_entry_valid_0; // @[TLB.scala 251:68]
  assign _GEN_359 = io_ptw_resp_bits_homogeneous ? _GEN_259 : superpage_entries_0_valid_0; // @[TLB.scala 251:68]
  assign _GEN_363 = io_ptw_resp_bits_homogeneous ? _GEN_263 : superpage_entries_1_valid_0; // @[TLB.scala 251:68]
  assign _GEN_367 = io_ptw_resp_bits_homogeneous ? _GEN_267 : superpage_entries_2_valid_0; // @[TLB.scala 251:68]
  assign _GEN_371 = io_ptw_resp_bits_homogeneous ? _GEN_271 : superpage_entries_3_valid_0; // @[TLB.scala 251:68]
  assign _GEN_373 = io_ptw_resp_bits_homogeneous ? _GEN_273 : sectored_entries_0_valid_0; // @[TLB.scala 251:68]
  assign _GEN_374 = io_ptw_resp_bits_homogeneous ? _GEN_274 : sectored_entries_0_valid_1; // @[TLB.scala 251:68]
  assign _GEN_375 = io_ptw_resp_bits_homogeneous ? _GEN_275 : sectored_entries_0_valid_2; // @[TLB.scala 251:68]
  assign _GEN_376 = io_ptw_resp_bits_homogeneous ? _GEN_276 : sectored_entries_0_valid_3; // @[TLB.scala 251:68]
  assign _GEN_383 = io_ptw_resp_bits_homogeneous ? _GEN_283 : sectored_entries_1_valid_0; // @[TLB.scala 251:68]
  assign _GEN_384 = io_ptw_resp_bits_homogeneous ? _GEN_284 : sectored_entries_1_valid_1; // @[TLB.scala 251:68]
  assign _GEN_385 = io_ptw_resp_bits_homogeneous ? _GEN_285 : sectored_entries_1_valid_2; // @[TLB.scala 251:68]
  assign _GEN_386 = io_ptw_resp_bits_homogeneous ? _GEN_286 : sectored_entries_1_valid_3; // @[TLB.scala 251:68]
  assign _GEN_393 = io_ptw_resp_bits_homogeneous ? _GEN_293 : sectored_entries_2_valid_0; // @[TLB.scala 251:68]
  assign _GEN_394 = io_ptw_resp_bits_homogeneous ? _GEN_294 : sectored_entries_2_valid_1; // @[TLB.scala 251:68]
  assign _GEN_395 = io_ptw_resp_bits_homogeneous ? _GEN_295 : sectored_entries_2_valid_2; // @[TLB.scala 251:68]
  assign _GEN_396 = io_ptw_resp_bits_homogeneous ? _GEN_296 : sectored_entries_2_valid_3; // @[TLB.scala 251:68]
  assign _GEN_403 = io_ptw_resp_bits_homogeneous ? _GEN_303 : sectored_entries_3_valid_0; // @[TLB.scala 251:68]
  assign _GEN_404 = io_ptw_resp_bits_homogeneous ? _GEN_304 : sectored_entries_3_valid_1; // @[TLB.scala 251:68]
  assign _GEN_405 = io_ptw_resp_bits_homogeneous ? _GEN_305 : sectored_entries_3_valid_2; // @[TLB.scala 251:68]
  assign _GEN_406 = io_ptw_resp_bits_homogeneous ? _GEN_306 : sectored_entries_3_valid_3; // @[TLB.scala 251:68]
  assign _GEN_413 = io_ptw_resp_bits_homogeneous ? _GEN_313 : sectored_entries_4_valid_0; // @[TLB.scala 251:68]
  assign _GEN_414 = io_ptw_resp_bits_homogeneous ? _GEN_314 : sectored_entries_4_valid_1; // @[TLB.scala 251:68]
  assign _GEN_415 = io_ptw_resp_bits_homogeneous ? _GEN_315 : sectored_entries_4_valid_2; // @[TLB.scala 251:68]
  assign _GEN_416 = io_ptw_resp_bits_homogeneous ? _GEN_316 : sectored_entries_4_valid_3; // @[TLB.scala 251:68]
  assign _GEN_423 = io_ptw_resp_bits_homogeneous ? _GEN_323 : sectored_entries_5_valid_0; // @[TLB.scala 251:68]
  assign _GEN_424 = io_ptw_resp_bits_homogeneous ? _GEN_324 : sectored_entries_5_valid_1; // @[TLB.scala 251:68]
  assign _GEN_425 = io_ptw_resp_bits_homogeneous ? _GEN_325 : sectored_entries_5_valid_2; // @[TLB.scala 251:68]
  assign _GEN_426 = io_ptw_resp_bits_homogeneous ? _GEN_326 : sectored_entries_5_valid_3; // @[TLB.scala 251:68]
  assign _GEN_433 = io_ptw_resp_bits_homogeneous ? _GEN_333 : sectored_entries_6_valid_0; // @[TLB.scala 251:68]
  assign _GEN_434 = io_ptw_resp_bits_homogeneous ? _GEN_334 : sectored_entries_6_valid_1; // @[TLB.scala 251:68]
  assign _GEN_435 = io_ptw_resp_bits_homogeneous ? _GEN_335 : sectored_entries_6_valid_2; // @[TLB.scala 251:68]
  assign _GEN_436 = io_ptw_resp_bits_homogeneous ? _GEN_336 : sectored_entries_6_valid_3; // @[TLB.scala 251:68]
  assign _GEN_443 = io_ptw_resp_bits_homogeneous ? _GEN_343 : sectored_entries_7_valid_0; // @[TLB.scala 251:68]
  assign _GEN_444 = io_ptw_resp_bits_homogeneous ? _GEN_344 : sectored_entries_7_valid_1; // @[TLB.scala 251:68]
  assign _GEN_445 = io_ptw_resp_bits_homogeneous ? _GEN_345 : sectored_entries_7_valid_2; // @[TLB.scala 251:68]
  assign _GEN_446 = io_ptw_resp_bits_homogeneous ? _GEN_346 : sectored_entries_7_valid_3; // @[TLB.scala 251:68]
  assign _GEN_455 = _T_1385 ? _GEN_355 : special_entry_valid_0; // @[TLB.scala 224:40]
  assign _GEN_459 = _T_1385 ? _GEN_359 : superpage_entries_0_valid_0; // @[TLB.scala 224:40]
  assign _GEN_463 = _T_1385 ? _GEN_363 : superpage_entries_1_valid_0; // @[TLB.scala 224:40]
  assign _GEN_467 = _T_1385 ? _GEN_367 : superpage_entries_2_valid_0; // @[TLB.scala 224:40]
  assign _GEN_471 = _T_1385 ? _GEN_371 : superpage_entries_3_valid_0; // @[TLB.scala 224:40]
  assign _GEN_473 = _T_1385 ? _GEN_373 : sectored_entries_0_valid_0; // @[TLB.scala 224:40]
  assign _GEN_474 = _T_1385 ? _GEN_374 : sectored_entries_0_valid_1; // @[TLB.scala 224:40]
  assign _GEN_475 = _T_1385 ? _GEN_375 : sectored_entries_0_valid_2; // @[TLB.scala 224:40]
  assign _GEN_476 = _T_1385 ? _GEN_376 : sectored_entries_0_valid_3; // @[TLB.scala 224:40]
  assign _GEN_483 = _T_1385 ? _GEN_383 : sectored_entries_1_valid_0; // @[TLB.scala 224:40]
  assign _GEN_484 = _T_1385 ? _GEN_384 : sectored_entries_1_valid_1; // @[TLB.scala 224:40]
  assign _GEN_485 = _T_1385 ? _GEN_385 : sectored_entries_1_valid_2; // @[TLB.scala 224:40]
  assign _GEN_486 = _T_1385 ? _GEN_386 : sectored_entries_1_valid_3; // @[TLB.scala 224:40]
  assign _GEN_493 = _T_1385 ? _GEN_393 : sectored_entries_2_valid_0; // @[TLB.scala 224:40]
  assign _GEN_494 = _T_1385 ? _GEN_394 : sectored_entries_2_valid_1; // @[TLB.scala 224:40]
  assign _GEN_495 = _T_1385 ? _GEN_395 : sectored_entries_2_valid_2; // @[TLB.scala 224:40]
  assign _GEN_496 = _T_1385 ? _GEN_396 : sectored_entries_2_valid_3; // @[TLB.scala 224:40]
  assign _GEN_503 = _T_1385 ? _GEN_403 : sectored_entries_3_valid_0; // @[TLB.scala 224:40]
  assign _GEN_504 = _T_1385 ? _GEN_404 : sectored_entries_3_valid_1; // @[TLB.scala 224:40]
  assign _GEN_505 = _T_1385 ? _GEN_405 : sectored_entries_3_valid_2; // @[TLB.scala 224:40]
  assign _GEN_506 = _T_1385 ? _GEN_406 : sectored_entries_3_valid_3; // @[TLB.scala 224:40]
  assign _GEN_513 = _T_1385 ? _GEN_413 : sectored_entries_4_valid_0; // @[TLB.scala 224:40]
  assign _GEN_514 = _T_1385 ? _GEN_414 : sectored_entries_4_valid_1; // @[TLB.scala 224:40]
  assign _GEN_515 = _T_1385 ? _GEN_415 : sectored_entries_4_valid_2; // @[TLB.scala 224:40]
  assign _GEN_516 = _T_1385 ? _GEN_416 : sectored_entries_4_valid_3; // @[TLB.scala 224:40]
  assign _GEN_523 = _T_1385 ? _GEN_423 : sectored_entries_5_valid_0; // @[TLB.scala 224:40]
  assign _GEN_524 = _T_1385 ? _GEN_424 : sectored_entries_5_valid_1; // @[TLB.scala 224:40]
  assign _GEN_525 = _T_1385 ? _GEN_425 : sectored_entries_5_valid_2; // @[TLB.scala 224:40]
  assign _GEN_526 = _T_1385 ? _GEN_426 : sectored_entries_5_valid_3; // @[TLB.scala 224:40]
  assign _GEN_533 = _T_1385 ? _GEN_433 : sectored_entries_6_valid_0; // @[TLB.scala 224:40]
  assign _GEN_534 = _T_1385 ? _GEN_434 : sectored_entries_6_valid_1; // @[TLB.scala 224:40]
  assign _GEN_535 = _T_1385 ? _GEN_435 : sectored_entries_6_valid_2; // @[TLB.scala 224:40]
  assign _GEN_536 = _T_1385 ? _GEN_436 : sectored_entries_6_valid_3; // @[TLB.scala 224:40]
  assign _GEN_543 = _T_1385 ? _GEN_443 : sectored_entries_7_valid_0; // @[TLB.scala 224:40]
  assign _GEN_544 = _T_1385 ? _GEN_444 : sectored_entries_7_valid_1; // @[TLB.scala 224:40]
  assign _GEN_545 = _T_1385 ? _GEN_445 : sectored_entries_7_valid_2; // @[TLB.scala 224:40]
  assign _GEN_546 = _T_1385 ? _GEN_446 : sectored_entries_7_valid_3; // @[TLB.scala 224:40]
  assign _T_2136 = {_GEN_55[11],_GEN_51[11],_GEN_47[11],_GEN_43[11],_GEN_39[11],_GEN_35[11]}; // @[Cat.scala 30:58]
  assign ptw_ae_array = {1'h0,special_entry_data_0[11],superpage_entries_3_data_0[11],superpage_entries_2_data_0[11],superpage_entries_1_data_0[11],superpage_entries_0_data_0[11],_GEN_63[11],_GEN_59[11],_T_2136}; // @[Cat.scala 30:58]
  assign _T_2145 = ~priv_s | io_ptw_status_sum; // @[TLB.scala 306:32]
  assign _T_2150 = {_GEN_55[13],_GEN_51[13],_GEN_47[13],_GEN_43[13],_GEN_39[13],_GEN_35[13]}; // @[Cat.scala 30:58]
  assign _T_2157 = {special_entry_data_0[13],superpage_entries_3_data_0[13],superpage_entries_2_data_0[13],superpage_entries_1_data_0[13],superpage_entries_0_data_0[13],_GEN_63[13],_GEN_59[13],_T_2150}; // @[Cat.scala 30:58]
  assign _T_2158 = _T_2145 ? _T_2157 : 13'h0; // @[TLB.scala 306:23]
  assign _T_2172 = priv_s ? ~_T_2157 : 13'h0; // @[TLB.scala 306:89]
  assign priv_rw_ok = _T_2158 | _T_2172; // @[TLB.scala 306:84]
  assign _T_2202 = {_GEN_55[8],_GEN_51[8],_GEN_47[8],_GEN_43[8],_GEN_39[8],_GEN_35[8]}; // @[Cat.scala 30:58]
  assign _T_2209 = {special_entry_data_0[8],superpage_entries_3_data_0[8],superpage_entries_2_data_0[8],superpage_entries_1_data_0[8],superpage_entries_0_data_0[8],_GEN_63[8],_GEN_59[8],_T_2202}; // @[Cat.scala 30:58]
  assign _T_2214 = {_GEN_55[9],_GEN_51[9],_GEN_47[9],_GEN_43[9],_GEN_39[9],_GEN_35[9]}; // @[Cat.scala 30:58]
  assign _T_2221 = {special_entry_data_0[9],superpage_entries_3_data_0[9],superpage_entries_2_data_0[9],superpage_entries_1_data_0[9],superpage_entries_0_data_0[9],_GEN_63[9],_GEN_59[9],_T_2214}; // @[Cat.scala 30:58]
  assign _T_2222 = io_ptw_status_mxr ? _T_2221 : 13'h0; // @[TLB.scala 308:73]
  assign _T_2223 = _T_2209 | _T_2222; // @[TLB.scala 308:68]
  assign _T_2224 = priv_rw_ok & _T_2223; // @[TLB.scala 308:40]
  assign r_array = {1'h1,_T_2224}; // @[Cat.scala 30:58]
  assign _T_2229 = {_GEN_55[10],_GEN_51[10],_GEN_47[10],_GEN_43[10],_GEN_39[10],_GEN_35[10]}; // @[Cat.scala 30:58]
  assign _T_2236 = {special_entry_data_0[10],superpage_entries_3_data_0[10],superpage_entries_2_data_0[10],superpage_entries_1_data_0[10],superpage_entries_0_data_0[10],_GEN_63[10],_GEN_59[10],_T_2229}; // @[Cat.scala 30:58]
  assign _T_2237 = priv_rw_ok & _T_2236; // @[TLB.scala 309:40]
  assign w_array = {1'h1,_T_2237}; // @[Cat.scala 30:58]
  assign _T_2252 = prot_r ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign _T_2257 = {_GEN_55[5],_GEN_51[5],_GEN_47[5],_GEN_43[5],_GEN_39[5],_GEN_35[5]}; // @[Cat.scala 30:58]
  assign _T_2264 = {_T_2252,superpage_entries_3_data_0[5],superpage_entries_2_data_0[5],superpage_entries_1_data_0[5],superpage_entries_0_data_0[5],_GEN_63[5],_GEN_59[5],_T_2257}; // @[Cat.scala 30:58]
  assign pr_array = _T_2264 | ptw_ae_array; // @[TLB.scala 311:87]
  assign _T_2266 = prot_w ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign _T_2271 = {_GEN_55[7],_GEN_51[7],_GEN_47[7],_GEN_43[7],_GEN_39[7],_GEN_35[7]}; // @[Cat.scala 30:58]
  assign _T_2278 = {_T_2266,superpage_entries_3_data_0[7],superpage_entries_2_data_0[7],superpage_entries_1_data_0[7],superpage_entries_0_data_0[7],_GEN_63[7],_GEN_59[7],_T_2271}; // @[Cat.scala 30:58]
  assign pw_array = _T_2278 | ptw_ae_array; // @[TLB.scala 312:87]
  assign _T_2294 = prot_al ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign _T_2299 = {_GEN_55[3],_GEN_51[3],_GEN_47[3],_GEN_43[3],_GEN_39[3],_GEN_35[3]}; // @[Cat.scala 30:58]
  assign paa_array = {_T_2294,superpage_entries_3_data_0[3],superpage_entries_2_data_0[3],superpage_entries_1_data_0[3],superpage_entries_0_data_0[3],_GEN_63[3],_GEN_59[3],_T_2299}; // @[Cat.scala 30:58]
  assign _T_2312 = {_GEN_55[4],_GEN_51[4],_GEN_47[4],_GEN_43[4],_GEN_39[4],_GEN_35[4]}; // @[Cat.scala 30:58]
  assign pal_array = {_T_2294,superpage_entries_3_data_0[4],superpage_entries_2_data_0[4],superpage_entries_1_data_0[4],superpage_entries_0_data_0[4],_GEN_63[4],_GEN_59[4],_T_2312}; // @[Cat.scala 30:58]
  assign _T_2320 = prot_eff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign _T_2325 = {_GEN_55[2],_GEN_51[2],_GEN_47[2],_GEN_43[2],_GEN_39[2],_GEN_35[2]}; // @[Cat.scala 30:58]
  assign eff_array = {_T_2320,superpage_entries_3_data_0[2],superpage_entries_2_data_0[2],superpage_entries_1_data_0[2],superpage_entries_0_data_0[2],_GEN_63[2],_GEN_59[2],_T_2325}; // @[Cat.scala 30:58]
  assign _T_2333 = cacheable ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign _T_2338 = {_GEN_55[1],_GEN_51[1],_GEN_47[1],_GEN_43[1],_GEN_39[1],_GEN_35[1]}; // @[Cat.scala 30:58]
  assign c_array = {_T_2333,superpage_entries_3_data_0[1],superpage_entries_2_data_0[1],superpage_entries_1_data_0[1],superpage_entries_0_data_0[1],_GEN_63[1],_GEN_59[1],_T_2338}; // @[Cat.scala 30:58]
  assign _T_2358 = 4'h1 << io_req_bits_size; // @[OneHot.scala 45:35]
  assign _T_2361 = _T_2358 - 4'h1; // @[TLB.scala 320:69]
  assign _GEN_1000 = {{36'd0}, _T_2361}; // @[TLB.scala 320:39]
  assign _T_2362 = io_req_bits_vaddr & _GEN_1000; // @[TLB.scala 320:39]
  assign misaligned = _T_2362 != 40'h0; // @[TLB.scala 320:75]
  assign _T_2364 = $signed(io_req_bits_vaddr) < 40'sh0; // @[TLB.scala 323:37]
  assign _T_2365 = io_req_bits_vaddr[38:12]; // @[TLB.scala 323:53]
  assign _T_2366 = $signed(_T_2365) < 27'sh0; // @[TLB.scala 323:60]
  assign _T_2367 = _T_2364 != _T_2366; // @[TLB.scala 323:44]
  assign bad_va = vm_enabled & _T_2367; // @[TLB.scala 321:27]
  assign _T_2368 = misaligned ? eff_array : 14'h0; // @[TLB.scala 327:8]
  assign _T_2369 = io_req_bits_cmd == 5'h6; // @[package.scala 14:47]
  assign _T_2370 = io_req_bits_cmd == 5'h7; // @[package.scala 14:47]
  assign _T_2371 = _T_2369 | _T_2370; // @[package.scala 14:62]
  assign _T_2374 = _T_2371 ? ~c_array : 14'h0; // @[TLB.scala 328:8]
  assign ae_array = _T_2368 | _T_2374; // @[TLB.scala 327:37]
  assign _T_2375 = io_req_bits_cmd == 5'h0; // @[Consts.scala 93:31]
  assign _T_2377 = _T_2375 | _T_2369; // @[Consts.scala 93:41]
  assign _T_2379 = _T_2377 | _T_2370; // @[Consts.scala 93:58]
  assign _T_2380 = io_req_bits_cmd == 5'h4; // @[package.scala 14:47]
  assign _T_2381 = io_req_bits_cmd == 5'h9; // @[package.scala 14:47]
  assign _T_2382 = io_req_bits_cmd == 5'ha; // @[package.scala 14:47]
  assign _T_2383 = io_req_bits_cmd == 5'hb; // @[package.scala 14:47]
  assign _T_2384 = _T_2380 | _T_2381; // @[package.scala 14:62]
  assign _T_2385 = _T_2384 | _T_2382; // @[package.scala 14:62]
  assign _T_2386 = _T_2385 | _T_2383; // @[package.scala 14:62]
  assign _T_2387 = io_req_bits_cmd == 5'h8; // @[package.scala 14:47]
  assign _T_2388 = io_req_bits_cmd == 5'hc; // @[package.scala 14:47]
  assign _T_2389 = io_req_bits_cmd == 5'hd; // @[package.scala 14:47]
  assign _T_2390 = io_req_bits_cmd == 5'he; // @[package.scala 14:47]
  assign _T_2391 = io_req_bits_cmd == 5'hf; // @[package.scala 14:47]
  assign _T_2392 = _T_2387 | _T_2388; // @[package.scala 14:62]
  assign _T_2393 = _T_2392 | _T_2389; // @[package.scala 14:62]
  assign _T_2394 = _T_2393 | _T_2390; // @[package.scala 14:62]
  assign _T_2395 = _T_2394 | _T_2391; // @[package.scala 14:62]
  assign _T_2396 = _T_2386 | _T_2395; // @[Consts.scala 91:44]
  assign _T_2397 = _T_2379 | _T_2396; // @[Consts.scala 93:75]
  assign _T_2399 = ae_array | ~pr_array; // @[TLB.scala 329:59]
  assign ae_ld_array = _T_2397 ? _T_2399 : 14'h0; // @[TLB.scala 329:24]
  assign _T_2400 = io_req_bits_cmd == 5'h1; // @[Consts.scala 94:32]
  assign _T_2401 = io_req_bits_cmd == 5'h11; // @[Consts.scala 94:49]
  assign _T_2402 = _T_2400 | _T_2401; // @[Consts.scala 94:42]
  assign _T_2404 = _T_2402 | _T_2370; // @[Consts.scala 94:59]
  assign _T_2422 = _T_2404 | _T_2396; // @[Consts.scala 94:76]
  assign _T_2424 = ae_array | ~pw_array; // @[TLB.scala 331:44]
  assign _T_2425 = _T_2422 ? _T_2424 : 14'h0; // @[TLB.scala 331:8]
  assign _T_2435 = _T_2386 ? ~pal_array : 14'h0; // @[TLB.scala 332:8]
  assign _T_2436 = _T_2425 | _T_2435; // @[TLB.scala 331:62]
  assign _T_2448 = _T_2395 ? ~paa_array : 14'h0; // @[TLB.scala 333:8]
  assign ae_st_array = _T_2436 | _T_2448; // @[TLB.scala 332:79]
  assign _T_2472 = misaligned & _T_2397; // @[TLB.scala 334:36]
  assign ma_ld_array = _T_2472 ? ~eff_array : 14'h0; // @[TLB.scala 334:24]
  assign _T_2497 = misaligned & _T_2422; // @[TLB.scala 335:36]
  assign ma_st_array = _T_2497 ? ~eff_array : 14'h0; // @[TLB.scala 335:24]
  assign _T_2522 = r_array | ptw_ae_array; // @[TLB.scala 336:60]
  assign pf_ld_array = _T_2397 ? ~_T_2522 : 14'h0; // @[TLB.scala 336:24]
  assign _T_2547 = w_array | ptw_ae_array; // @[TLB.scala 337:61]
  assign pf_st_array = _T_2422 ? ~_T_2547 : 14'h0; // @[TLB.scala 337:24]
  assign tlb_hit = real_hits != 13'h0; // @[TLB.scala 340:27]
  assign _T_2551 = vm_enabled & ~bad_va; // @[TLB.scala 341:29]
  assign tlb_miss = _T_2551 & ~tlb_hit; // @[TLB.scala 341:40]
  assign _T_2557 = io_req_valid & vm_enabled; // @[TLB.scala 345:22]
  assign _T_2558 = sector_hits_0 | sector_hits_1; // @[package.scala 63:59]
  assign _T_2559 = _T_2558 | sector_hits_2; // @[package.scala 63:59]
  assign _T_2560 = _T_2559 | sector_hits_3; // @[package.scala 63:59]
  assign _T_2561 = _T_2560 | sector_hits_4; // @[package.scala 63:59]
  assign _T_2562 = _T_2561 | sector_hits_5; // @[package.scala 63:59]
  assign _T_2563 = _T_2562 | sector_hits_6; // @[package.scala 63:59]
  assign _T_2564 = _T_2563 | sector_hits_7; // @[package.scala 63:59]
  assign _T_2571 = {sector_hits_7,sector_hits_6,sector_hits_5,sector_hits_4,sector_hits_3,sector_hits_2,sector_hits_1,sector_hits_0}; // @[Cat.scala 30:58]
  assign _T_2574 = _T_2571[7:4] != 4'h0; // @[OneHot.scala 28:14]
  assign _T_2575 = _T_2571[7:4] | _T_2571[3:0]; // @[OneHot.scala 28:28]
  assign _T_2578 = _T_2575[3:2] != 2'h0; // @[OneHot.scala 28:14]
  assign _T_2579 = _T_2575[3:2] | _T_2575[1:0]; // @[OneHot.scala 28:28]
  assign _T_2582 = {_T_2574,_T_2578,_T_2579[1]}; // @[Cat.scala 30:58]
  assign _T_2583 = {_T_2554, 1'h0}; // @[Replacement.scala 46:28]
  assign _T_2587 = _T_2583 | 8'h2; // @[Replacement.scala 50:37]
  assign _T_2589 = ~_T_2583 | 8'h2; // @[Replacement.scala 50:37]
  assign _T_2591 = _T_2582[2] ? ~_T_2589 : _T_2587; // @[Replacement.scala 50:37]
  assign _T_2592 = {1'h1,_T_2582[2]}; // @[Cat.scala 30:58]
  assign _T_2595 = 4'h1 << _T_2592; // @[Replacement.scala 50:37]
  assign _GEN_1001 = {{4'd0}, _T_2595}; // @[Replacement.scala 50:37]
  assign _T_2596 = _T_2591 | _GEN_1001; // @[Replacement.scala 50:37]
  assign _T_2598 = ~_T_2591 | _GEN_1001; // @[Replacement.scala 50:37]
  assign _T_2600 = _T_2582[1] ? ~_T_2598 : _T_2596; // @[Replacement.scala 50:37]
  assign _T_2601 = {1'h1,_T_2582[2],_T_2582[1]}; // @[Cat.scala 30:58]
  assign _T_2604 = 8'h1 << _T_2601; // @[Replacement.scala 50:37]
  assign _T_2605 = _T_2600 | _T_2604; // @[Replacement.scala 50:37]
  assign _T_2607 = ~_T_2600 | _T_2604; // @[Replacement.scala 50:37]
  assign _T_2609 = _T_2582[0] ? ~_T_2607 : _T_2605; // @[Replacement.scala 50:37]
  assign _T_2612 = superpage_hits_0 | superpage_hits_1; // @[package.scala 63:59]
  assign _T_2613 = _T_2612 | superpage_hits_2; // @[package.scala 63:59]
  assign _T_2614 = _T_2613 | superpage_hits_3; // @[package.scala 63:59]
  assign _T_2617 = {superpage_hits_3,superpage_hits_2,superpage_hits_1,superpage_hits_0}; // @[Cat.scala 30:58]
  assign _T_2620 = _T_2617[3:2] != 2'h0; // @[OneHot.scala 28:14]
  assign _T_2621 = _T_2617[3:2] | _T_2617[1:0]; // @[OneHot.scala 28:28]
  assign _T_2623 = {_T_2620,_T_2621[1]}; // @[Cat.scala 30:58]
  assign _T_2624 = {_T_2556, 1'h0}; // @[Replacement.scala 46:28]
  assign _T_2628 = _T_2624 | 4'h2; // @[Replacement.scala 50:37]
  assign _T_2630 = ~_T_2624 | 4'h2; // @[Replacement.scala 50:37]
  assign _T_2632 = _T_2623[1] ? ~_T_2630 : _T_2628; // @[Replacement.scala 50:37]
  assign _T_2633 = {1'h1,_T_2623[1]}; // @[Cat.scala 30:58]
  assign _T_2636 = 4'h1 << _T_2633; // @[Replacement.scala 50:37]
  assign _T_2637 = _T_2632 | _T_2636; // @[Replacement.scala 50:37]
  assign _T_2639 = ~_T_2632 | _T_2636; // @[Replacement.scala 50:37]
  assign _T_2641 = _T_2623[0] ? ~_T_2639 : _T_2637; // @[Replacement.scala 50:37]
  assign _T_2653 = real_hits[1] | real_hits[2]; // @[Misc.scala 187:16]
  assign _T_2655 = real_hits[1] & real_hits[2]; // @[Misc.scala 187:61]
  assign _T_2657 = real_hits[0] | _T_2653; // @[Misc.scala 187:16]
  assign _T_2659 = real_hits[0] & _T_2653; // @[Misc.scala 187:61]
  assign _T_2660 = _T_2655 | _T_2659; // @[Misc.scala 187:49]
  assign _T_2669 = real_hits[4] | real_hits[5]; // @[Misc.scala 187:16]
  assign _T_2671 = real_hits[4] & real_hits[5]; // @[Misc.scala 187:61]
  assign _T_2673 = real_hits[3] | _T_2669; // @[Misc.scala 187:16]
  assign _T_2675 = real_hits[3] & _T_2669; // @[Misc.scala 187:61]
  assign _T_2676 = _T_2671 | _T_2675; // @[Misc.scala 187:49]
  assign _T_2677 = _T_2657 | _T_2673; // @[Misc.scala 187:16]
  assign _T_2678 = _T_2660 | _T_2676; // @[Misc.scala 187:37]
  assign _T_2679 = _T_2657 & _T_2673; // @[Misc.scala 187:61]
  assign _T_2680 = _T_2678 | _T_2679; // @[Misc.scala 187:49]
  assign _T_2690 = real_hits[7] | real_hits[8]; // @[Misc.scala 187:16]
  assign _T_2692 = real_hits[7] & real_hits[8]; // @[Misc.scala 187:61]
  assign _T_2694 = real_hits[6] | _T_2690; // @[Misc.scala 187:16]
  assign _T_2696 = real_hits[6] & _T_2690; // @[Misc.scala 187:61]
  assign _T_2697 = _T_2692 | _T_2696; // @[Misc.scala 187:49]
  assign _T_2704 = real_hits[9] | real_hits[10]; // @[Misc.scala 187:16]
  assign _T_2706 = real_hits[9] & real_hits[10]; // @[Misc.scala 187:61]
  assign _T_2713 = real_hits[11] | real_hits[12]; // @[Misc.scala 187:16]
  assign _T_2715 = real_hits[11] & real_hits[12]; // @[Misc.scala 187:61]
  assign _T_2717 = _T_2704 | _T_2713; // @[Misc.scala 187:16]
  assign _T_2718 = _T_2706 | _T_2715; // @[Misc.scala 187:37]
  assign _T_2719 = _T_2704 & _T_2713; // @[Misc.scala 187:61]
  assign _T_2720 = _T_2718 | _T_2719; // @[Misc.scala 187:49]
  assign _T_2721 = _T_2694 | _T_2717; // @[Misc.scala 187:16]
  assign _T_2722 = _T_2697 | _T_2720; // @[Misc.scala 187:37]
  assign _T_2723 = _T_2694 & _T_2717; // @[Misc.scala 187:61]
  assign _T_2724 = _T_2722 | _T_2723; // @[Misc.scala 187:49]
  assign _T_2726 = _T_2680 | _T_2724; // @[Misc.scala 187:37]
  assign _T_2727 = _T_2677 & _T_2721; // @[Misc.scala 187:61]
  assign multipleHits = _T_2726 | _T_2727; // @[Misc.scala 187:49]
  assign _T_2752 = bad_va & _T_2397; // @[TLB.scala 358:28]
  assign _T_2753 = pf_ld_array & hits; // @[TLB.scala 358:72]
  assign _T_2754 = _T_2753 != 14'h0; // @[TLB.scala 358:80]
  assign _T_2779 = bad_va & _T_2422; // @[TLB.scala 359:28]
  assign _T_2780 = pf_st_array & hits; // @[TLB.scala 359:73]
  assign _T_2781 = _T_2780 != 14'h0; // @[TLB.scala 359:81]
  assign _T_2786 = ae_ld_array & hits; // @[TLB.scala 361:33]
  assign _T_2788 = ae_st_array & hits; // @[TLB.scala 362:33]
  assign _T_2793 = ma_ld_array & hits; // @[TLB.scala 364:33]
  assign _T_2795 = ma_st_array & hits; // @[TLB.scala 365:33]
  assign _T_2797 = c_array & hits; // @[TLB.scala 367:33]
  assign _T_2802 = io_ptw_resp_valid | tlb_miss; // @[TLB.scala 369:29]
  assign _T_2808 = io_req_ready & io_req_valid; // @[Decoupled.scala 37:37]
  assign _T_2809 = _T_2808 & tlb_miss; // @[TLB.scala 385:25]
  assign _T_2814 = {{1'd0}, _T_2624[3:1]}; // @[Replacement.scala 61:48]
  assign _T_2817 = {1'h1,_T_2814[0]}; // @[Cat.scala 30:58]
  assign _T_2821 = _T_2624 >> _T_2817; // @[Replacement.scala 61:48]
  assign _T_2824 = {1'h1,_T_2814[0],_T_2821[0]}; // @[Cat.scala 30:58]
  assign _T_2828 = {superpage_entries_3_valid_0,superpage_entries_2_valid_0,superpage_entries_1_valid_0,superpage_entries_0_valid_0}; // @[Cat.scala 30:58]
  assign _T_2830 = ~_T_2828 == 4'h0; // @[TLB.scala 440:16]
  assign _T_2832 = ~_T_2828[0]; // @[OneHot.scala 39:40]
  assign _T_2833 = ~_T_2828[1]; // @[OneHot.scala 39:40]
  assign _T_2834 = ~_T_2828[2]; // @[OneHot.scala 39:40]
  assign _T_2844 = {{1'd0}, _T_2583[7:1]}; // @[Replacement.scala 61:48]
  assign _T_2847 = {1'h1,_T_2844[0]}; // @[Cat.scala 30:58]
  assign _T_2851 = _T_2583 >> _T_2847; // @[Replacement.scala 61:48]
  assign _T_2854 = {1'h1,_T_2844[0],_T_2851[0]}; // @[Cat.scala 30:58]
  assign _T_2858 = _T_2583 >> _T_2854; // @[Replacement.scala 61:48]
  assign _T_2861 = {1'h1,_T_2844[0],_T_2851[0],_T_2858[0]}; // @[Cat.scala 30:58]
  assign _T_2893 = {_T_766,_T_760,_T_754,_T_748,_T_742,_T_736,_T_730,_T_724}; // @[Cat.scala 30:58]
  assign _T_2895 = ~_T_2893 == 8'h0; // @[TLB.scala 440:16]
  assign _T_2897 = ~_T_2893[0]; // @[OneHot.scala 39:40]
  assign _T_2898 = ~_T_2893[1]; // @[OneHot.scala 39:40]
  assign _T_2899 = ~_T_2893[2]; // @[OneHot.scala 39:40]
  assign _T_2900 = ~_T_2893[3]; // @[OneHot.scala 39:40]
  assign _T_2901 = ~_T_2893[4]; // @[OneHot.scala 39:40]
  assign _T_2902 = ~_T_2893[5]; // @[OneHot.scala 39:40]
  assign _T_2903 = ~_T_2893[6]; // @[OneHot.scala 39:40]
  assign _T_2940 = state == 2'h2; // @[TLB.scala 399:17]
  assign _T_2941 = _T_2940 & io_sfence_valid; // @[TLB.scala 399:28]
  assign _T_2946 = io_sfence_bits_addr[38:12] == vpn; // @[TLB.scala 414:72]
  assign _T_2947 = ~io_sfence_bits_rs1 | _T_2946; // @[TLB.scala 414:34]
  assign _T_2949 = _T_2947 | reset; // @[TLB.scala 414:13]
  assign _T_2957 = _T_725[26:18] == 9'h0; // @[TLB.scala 150:63]
  assign _GEN_652 = sectored_entries_0_data_0[12] ? _GEN_473 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_653 = sectored_entries_0_data_1[12] ? _GEN_474 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_654 = sectored_entries_0_data_2[12] ? _GEN_475 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_655 = sectored_entries_0_data_3[12] ? _GEN_476 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_656 = io_sfence_bits_rs2 & _GEN_652; // @[TLB.scala 417:40]
  assign _GEN_657 = io_sfence_bits_rs2 & _GEN_653; // @[TLB.scala 417:40]
  assign _GEN_658 = io_sfence_bits_rs2 & _GEN_654; // @[TLB.scala 417:40]
  assign _GEN_659 = io_sfence_bits_rs2 & _GEN_655; // @[TLB.scala 417:40]
  assign _T_3128 = _T_731[26:18] == 9'h0; // @[TLB.scala 150:63]
  assign _GEN_680 = sectored_entries_1_data_0[12] ? _GEN_483 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_681 = sectored_entries_1_data_1[12] ? _GEN_484 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_682 = sectored_entries_1_data_2[12] ? _GEN_485 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_683 = sectored_entries_1_data_3[12] ? _GEN_486 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_684 = io_sfence_bits_rs2 & _GEN_680; // @[TLB.scala 417:40]
  assign _GEN_685 = io_sfence_bits_rs2 & _GEN_681; // @[TLB.scala 417:40]
  assign _GEN_686 = io_sfence_bits_rs2 & _GEN_682; // @[TLB.scala 417:40]
  assign _GEN_687 = io_sfence_bits_rs2 & _GEN_683; // @[TLB.scala 417:40]
  assign _T_3299 = _T_737[26:18] == 9'h0; // @[TLB.scala 150:63]
  assign _GEN_708 = sectored_entries_2_data_0[12] ? _GEN_493 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_709 = sectored_entries_2_data_1[12] ? _GEN_494 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_710 = sectored_entries_2_data_2[12] ? _GEN_495 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_711 = sectored_entries_2_data_3[12] ? _GEN_496 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_712 = io_sfence_bits_rs2 & _GEN_708; // @[TLB.scala 417:40]
  assign _GEN_713 = io_sfence_bits_rs2 & _GEN_709; // @[TLB.scala 417:40]
  assign _GEN_714 = io_sfence_bits_rs2 & _GEN_710; // @[TLB.scala 417:40]
  assign _GEN_715 = io_sfence_bits_rs2 & _GEN_711; // @[TLB.scala 417:40]
  assign _T_3470 = _T_743[26:18] == 9'h0; // @[TLB.scala 150:63]
  assign _GEN_736 = sectored_entries_3_data_0[12] ? _GEN_503 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_737 = sectored_entries_3_data_1[12] ? _GEN_504 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_738 = sectored_entries_3_data_2[12] ? _GEN_505 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_739 = sectored_entries_3_data_3[12] ? _GEN_506 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_740 = io_sfence_bits_rs2 & _GEN_736; // @[TLB.scala 417:40]
  assign _GEN_741 = io_sfence_bits_rs2 & _GEN_737; // @[TLB.scala 417:40]
  assign _GEN_742 = io_sfence_bits_rs2 & _GEN_738; // @[TLB.scala 417:40]
  assign _GEN_743 = io_sfence_bits_rs2 & _GEN_739; // @[TLB.scala 417:40]
  assign _T_3641 = _T_749[26:18] == 9'h0; // @[TLB.scala 150:63]
  assign _GEN_764 = sectored_entries_4_data_0[12] ? _GEN_513 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_765 = sectored_entries_4_data_1[12] ? _GEN_514 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_766 = sectored_entries_4_data_2[12] ? _GEN_515 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_767 = sectored_entries_4_data_3[12] ? _GEN_516 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_768 = io_sfence_bits_rs2 & _GEN_764; // @[TLB.scala 417:40]
  assign _GEN_769 = io_sfence_bits_rs2 & _GEN_765; // @[TLB.scala 417:40]
  assign _GEN_770 = io_sfence_bits_rs2 & _GEN_766; // @[TLB.scala 417:40]
  assign _GEN_771 = io_sfence_bits_rs2 & _GEN_767; // @[TLB.scala 417:40]
  assign _T_3812 = _T_755[26:18] == 9'h0; // @[TLB.scala 150:63]
  assign _GEN_792 = sectored_entries_5_data_0[12] ? _GEN_523 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_793 = sectored_entries_5_data_1[12] ? _GEN_524 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_794 = sectored_entries_5_data_2[12] ? _GEN_525 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_795 = sectored_entries_5_data_3[12] ? _GEN_526 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_796 = io_sfence_bits_rs2 & _GEN_792; // @[TLB.scala 417:40]
  assign _GEN_797 = io_sfence_bits_rs2 & _GEN_793; // @[TLB.scala 417:40]
  assign _GEN_798 = io_sfence_bits_rs2 & _GEN_794; // @[TLB.scala 417:40]
  assign _GEN_799 = io_sfence_bits_rs2 & _GEN_795; // @[TLB.scala 417:40]
  assign _T_3983 = _T_761[26:18] == 9'h0; // @[TLB.scala 150:63]
  assign _GEN_820 = sectored_entries_6_data_0[12] ? _GEN_533 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_821 = sectored_entries_6_data_1[12] ? _GEN_534 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_822 = sectored_entries_6_data_2[12] ? _GEN_535 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_823 = sectored_entries_6_data_3[12] ? _GEN_536 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_824 = io_sfence_bits_rs2 & _GEN_820; // @[TLB.scala 417:40]
  assign _GEN_825 = io_sfence_bits_rs2 & _GEN_821; // @[TLB.scala 417:40]
  assign _GEN_826 = io_sfence_bits_rs2 & _GEN_822; // @[TLB.scala 417:40]
  assign _GEN_827 = io_sfence_bits_rs2 & _GEN_823; // @[TLB.scala 417:40]
  assign _T_4154 = _T_767[26:18] == 9'h0; // @[TLB.scala 150:63]
  assign _GEN_848 = sectored_entries_7_data_0[12] ? _GEN_543 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_849 = sectored_entries_7_data_1[12] ? _GEN_544 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_850 = sectored_entries_7_data_2[12] ? _GEN_545 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_851 = sectored_entries_7_data_3[12] ? _GEN_546 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_852 = io_sfence_bits_rs2 & _GEN_848; // @[TLB.scala 417:40]
  assign _GEN_853 = io_sfence_bits_rs2 & _GEN_849; // @[TLB.scala 417:40]
  assign _GEN_854 = io_sfence_bits_rs2 & _GEN_850; // @[TLB.scala 417:40]
  assign _GEN_855 = io_sfence_bits_rs2 & _GEN_851; // @[TLB.scala 417:40]
  assign _GEN_861 = superpage_entries_0_data_0[12] ? _GEN_459 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_862 = io_sfence_bits_rs2 & _GEN_861; // @[TLB.scala 417:40]
  assign _GEN_865 = superpage_entries_1_data_0[12] ? _GEN_463 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_866 = io_sfence_bits_rs2 & _GEN_865; // @[TLB.scala 417:40]
  assign _GEN_869 = superpage_entries_2_data_0[12] ? _GEN_467 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_870 = io_sfence_bits_rs2 & _GEN_869; // @[TLB.scala 417:40]
  assign _GEN_873 = superpage_entries_3_data_0[12] ? _GEN_471 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_874 = io_sfence_bits_rs2 & _GEN_873; // @[TLB.scala 417:40]
  assign _GEN_877 = special_entry_data_0[12] ? _GEN_455 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_878 = io_sfence_bits_rs2 & _GEN_877; // @[TLB.scala 417:40]
  assign _T_4530 = multipleHits | reset; // @[TLB.scala 421:24]
  assign io_req_ready = state == 2'h0; // @[TLB.scala 357:16]
  assign io_resp_miss = _T_2802 | multipleHits; // @[TLB.scala 369:16]
  assign io_resp_paddr = {ppn,io_req_bits_vaddr[11:0]}; // @[TLB.scala 370:17]
  assign io_resp_pf_ld = _T_2752 | _T_2754; // @[TLB.scala 358:17]
  assign io_resp_pf_st = _T_2779 | _T_2781; // @[TLB.scala 359:17]
  assign io_resp_ae_ld = _T_2786 != 14'h0; // @[TLB.scala 361:17]
  assign io_resp_ae_st = _T_2788 != 14'h0; // @[TLB.scala 362:17]
  assign io_resp_ma_ld = _T_2793 != 14'h0; // @[TLB.scala 364:17]
  assign io_resp_ma_st = _T_2795 != 14'h0; // @[TLB.scala 365:17]
  assign io_resp_cacheable = _T_2797 != 14'h0; // @[TLB.scala 367:21]
  assign io_ptw_req_valid = state == 2'h1; // @[TLB.scala 372:20]
  assign io_ptw_req_bits_valid = 1'h1; // @[TLB.scala 373:25]
  assign io_ptw_req_bits_bits_addr = r_refill_tag; // @[TLB.scala 374:29]
  assign pmp_io_prv = _T_363 ? 2'h1 : io_ptw_status_dprv; // @[TLB.scala 194:14]
  assign pmp_io_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_addr = io_ptw_pmp_0_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_mask = io_ptw_pmp_0_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_addr = io_ptw_pmp_1_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_mask = io_ptw_pmp_1_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_addr = io_ptw_pmp_2_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_mask = io_ptw_pmp_2_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_addr = io_ptw_pmp_3_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_mask = io_ptw_pmp_3_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_addr = io_ptw_pmp_4_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_mask = io_ptw_pmp_4_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_addr = io_ptw_pmp_5_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_mask = io_ptw_pmp_5_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_addr = io_ptw_pmp_6_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_mask = io_ptw_pmp_6_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_addr = io_ptw_pmp_7_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_mask = io_ptw_pmp_7_mask; // @[TLB.scala 193:14]
  assign pmp_io_addr = mpu_physaddr[31:0]; // @[TLB.scala 191:15]
  assign pmp_io_size = io_req_bits_size; // @[TLB.scala 192:15]
  assign TLB_cov_read_addr = TLB_state;
  assign TLB_cov_read_data = TLB_cov[TLB_cov_read_addr]; // @[Coverage map for TLB]
  assign TLB_cov_write_data = 1'h1;
  assign TLB_cov_write_addr = TLB_state;
  assign TLB_cov_write_mask = 1'h1;
  assign TLB_cov_write_en = 1'h1;
  assign mux_cond_0 = sectored_entries_0_data_0[0];
  assign mux_cond_1 = ~sectored_entries_3_data_3[12];
  assign mux_cond_2 = prot_eff;
  assign mux_cond_3 = sectored_entries_1_data_0[0];
  assign mux_cond_4 = ~sectored_entries_4_data_3[12];
  assign mux_cond_5 = ~superpage_entries_0_data_0[12];
  assign mux_cond_6 = ~sectored_entries_2_data_1[12];
  assign mux_cond_7 = sectored_entries_2_data_3[0];
  assign mux_cond_8 = prot_r;
  assign mux_cond_9 = ~sectored_entries_4_data_2[12];
  assign mux_cond_10 = ~sectored_entries_5_data_1[12];
  assign mux_cond_11 = sectored_entries_0_data_1[0];
  assign mux_cond_12 = sectored_entries_3_data_1[0];
  assign mux_cond_13 = ~sectored_entries_4_data_1[12];
  assign mux_cond_14 = sectored_entries_7_data_1[0];
  assign mux_cond_15 = ~sectored_entries_0_data_3[12];
  assign mux_cond_16 = ~sectored_entries_1_data_2[12];
  assign mux_cond_17 = sectored_entries_5_data_2[0];
  assign mux_cond_18 = ~special_entry_data_0[12];
  assign mux_cond_19 = sectored_entries_5_data_3[0];
  assign mux_cond_20 = sectored_entries_6_data_1[0];
  assign mux_cond_21 = ~sectored_entries_2_data_3[12];
  assign mux_cond_22 = ~superpage_entries_1_data_0[12];
  assign mux_cond_23 = ~sectored_entries_3_data_0[12];
  assign mux_cond_24 = sectored_entries_4_data_0[0];
  assign mux_cond_25 = sectored_entries_7_data_3[0];
  assign mux_cond_26 = ~sectored_entries_1_data_1[12];
  assign mux_cond_27 = sectored_entries_2_data_0[0];
  assign mux_cond_28 = ~sectored_entries_1_data_0[12];
  assign mux_cond_29 = sectored_entries_1_data_2[0];
  assign mux_cond_30 = ~sectored_entries_5_data_2[12];
  assign mux_cond_31 = sectored_entries_3_data_2[0];
  assign mux_cond_32 = ~sectored_entries_3_data_2[12];
  assign mux_cond_33 = ~sectored_entries_7_data_2[12];
  assign mux_cond_34 = ~sectored_entries_2_data_2[12];
  assign mux_cond_35 = sectored_entries_4_data_3[0];
  assign mux_cond_36 = sectored_entries_5_data_0[0];
  assign mux_cond_37 = sectored_entries_7_data_0[0];
  assign mux_cond_38 = sectored_entries_2_data_2[0];
  assign mux_cond_39 = sectored_entries_6_data_3[0];
  assign mux_cond_40 = ~superpage_entries_3_data_0[12];
  assign mux_cond_41 = ~sectored_entries_7_data_3[12];
  assign mux_cond_42 = ~sectored_entries_7_data_1[12];
  assign mux_cond_43 = sectored_entries_1_data_1[0];
  assign mux_cond_44 = prot_w;
  assign mux_cond_45 = sectored_entries_0_data_3[0];
  assign mux_cond_46 = cacheable;
  assign mux_cond_47 = sectored_entries_5_data_1[0];
  assign mux_cond_48 = ~sectored_entries_5_data_3[12];
  assign mux_cond_49 = ~sectored_entries_0_data_2[12];
  assign mux_cond_50 = ~sectored_entries_1_data_3[12];
  assign mux_cond_51 = sectored_entries_6_data_2[0];
  assign mux_cond_52 = ~sectored_entries_4_data_0[12];
  assign mux_cond_53 = ~sectored_entries_0_data_0[12];
  assign mux_cond_54 = ~sectored_entries_7_data_0[12];
  assign mux_cond_55 = ~sectored_entries_3_data_1[12];
  assign mux_cond_56 = ~sectored_entries_5_data_0[12];
  assign mux_cond_57 = sectored_entries_3_data_0[0];
  assign mux_cond_58 = sectored_entries_7_data_2[0];
  assign mux_cond_59 = ~sectored_entries_2_data_0[12];
  assign mux_cond_60 = sectored_entries_4_data_2[0];
  assign mux_cond_61 = sectored_entries_1_data_3[0];
  assign mux_cond_62 = ~sectored_entries_6_data_2[12];
  assign mux_cond_63 = ~sectored_entries_6_data_0[12];
  assign mux_cond_64 = ~sectored_entries_0_data_1[12];
  assign mux_cond_65 = sectored_entries_3_data_3[0];
  assign mux_cond_66 = ~superpage_entries_2_data_0[12];
  assign mux_cond_67 = sectored_entries_6_data_0[0];
  assign mux_cond_68 = sectored_entries_4_data_1[0];
  assign mux_cond_69 = ~sectored_entries_6_data_3[12];
  assign mux_cond_70 = sectored_entries_0_data_2[0];
  assign mux_cond_71 = sectored_entries_2_data_1[0];
  assign mux_cond_72 = ~sectored_entries_6_data_1[12];
  assign mux_cond_73 = prot_al;
  assign r_superpage_repl_addr_shl = {r_superpage_repl_addr, 8'h0};
  assign r_superpage_repl_addr_pad = {10'h0,r_superpage_repl_addr_shl};
  assign state_shl = {state, 1'h0};
  assign state_pad = {17'h0,state_shl};
  assign r_sectored_repl_addr_shl = {r_sectored_repl_addr, 13'h0};
  assign r_sectored_repl_addr_pad = {4'h0,r_sectored_repl_addr_shl};
  assign r_sectored_hit_addr_shl = {r_sectored_hit_addr, 5'h0};
  assign r_sectored_hit_addr_pad = {12'h0,r_sectored_hit_addr_shl};
  assign special_entry_valid_0_shl = {special_entry_valid_0, 10'h0};
  assign special_entry_valid_0_pad = {9'h0,special_entry_valid_0_shl};
  assign special_entry_level_shl = special_entry_level;
  assign special_entry_level_pad = {18'h0,special_entry_level_shl};
  assign r_sectored_hit_shl = {r_sectored_hit, 19'h0};
  assign r_sectored_hit_pad = r_sectored_hit_shl;
  assign mux_cond_0_shl = {mux_cond_0, 9'h0};
  assign mux_cond_0_pad = {10'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 18'h0};
  assign mux_cond_1_pad = {1'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 4'h0};
  assign mux_cond_2_pad = {15'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 5'h0};
  assign mux_cond_3_pad = {14'h0,mux_cond_3_shl};
  assign mux_cond_4_shl = {mux_cond_4, 15'h0};
  assign mux_cond_4_pad = {4'h0,mux_cond_4_shl};
  assign mux_cond_5_shl = {mux_cond_5, 2'h0};
  assign mux_cond_5_pad = {17'h0,mux_cond_5_shl};
  assign mux_cond_6_shl = {mux_cond_6, 1'h0};
  assign mux_cond_6_pad = {18'h0,mux_cond_6_shl};
  assign mux_cond_7_shl = {mux_cond_7, 9'h0};
  assign mux_cond_7_pad = {10'h0,mux_cond_7_shl};
  assign mux_cond_8_shl = {mux_cond_8, 5'h0};
  assign mux_cond_8_pad = {14'h0,mux_cond_8_shl};
  assign mux_cond_9_shl = {mux_cond_9, 5'h0};
  assign mux_cond_9_pad = {14'h0,mux_cond_9_shl};
  assign mux_cond_10_shl = {mux_cond_10, 7'h0};
  assign mux_cond_10_pad = {12'h0,mux_cond_10_shl};
  assign mux_cond_11_shl = {mux_cond_11, 1'h0};
  assign mux_cond_11_pad = {18'h0,mux_cond_11_shl};
  assign mux_cond_12_shl = {mux_cond_12, 14'h0};
  assign mux_cond_12_pad = {5'h0,mux_cond_12_shl};
  assign mux_cond_13_shl = {mux_cond_13, 11'h0};
  assign mux_cond_13_pad = {8'h0,mux_cond_13_shl};
  assign mux_cond_14_shl = {mux_cond_14, 2'h0};
  assign mux_cond_14_pad = {17'h0,mux_cond_14_shl};
  assign mux_cond_15_shl = {mux_cond_15, 17'h0};
  assign mux_cond_15_pad = {2'h0,mux_cond_15_shl};
  assign mux_cond_16_shl = mux_cond_16;
  assign mux_cond_16_pad = {19'h0,mux_cond_16_shl};
  assign mux_cond_17_shl = {mux_cond_17, 18'h0};
  assign mux_cond_17_pad = {1'h0,mux_cond_17_shl};
  assign mux_cond_18_shl = {mux_cond_18, 19'h0};
  assign mux_cond_18_pad = mux_cond_18_shl;
  assign mux_cond_19_shl = {mux_cond_19, 8'h0};
  assign mux_cond_19_pad = {11'h0,mux_cond_19_shl};
  assign mux_cond_20_shl = {mux_cond_20, 17'h0};
  assign mux_cond_20_pad = {2'h0,mux_cond_20_shl};
  assign mux_cond_21_shl = {mux_cond_21, 3'h0};
  assign mux_cond_21_pad = {16'h0,mux_cond_21_shl};
  assign mux_cond_22_shl = {mux_cond_22, 5'h0};
  assign mux_cond_22_pad = {14'h0,mux_cond_22_shl};
  assign mux_cond_23_shl = {mux_cond_23, 5'h0};
  assign mux_cond_23_pad = {14'h0,mux_cond_23_shl};
  assign mux_cond_24_shl = {mux_cond_24, 15'h0};
  assign mux_cond_24_pad = {4'h0,mux_cond_24_shl};
  assign mux_cond_25_shl = {mux_cond_25, 18'h0};
  assign mux_cond_25_pad = {1'h0,mux_cond_25_shl};
  assign mux_cond_26_shl = {mux_cond_26, 3'h0};
  assign mux_cond_26_pad = {16'h0,mux_cond_26_shl};
  assign mux_cond_27_shl = {mux_cond_27, 12'h0};
  assign mux_cond_27_pad = {7'h0,mux_cond_27_shl};
  assign mux_cond_28_shl = {mux_cond_28, 10'h0};
  assign mux_cond_28_pad = {9'h0,mux_cond_28_shl};
  assign mux_cond_29_shl = {mux_cond_29, 3'h0};
  assign mux_cond_29_pad = {16'h0,mux_cond_29_shl};
  assign mux_cond_30_shl = mux_cond_30;
  assign mux_cond_30_pad = {19'h0,mux_cond_30_shl};
  assign mux_cond_31_shl = {mux_cond_31, 18'h0};
  assign mux_cond_31_pad = {1'h0,mux_cond_31_shl};
  assign mux_cond_32_shl = {mux_cond_32, 12'h0};
  assign mux_cond_32_pad = {7'h0,mux_cond_32_shl};
  assign mux_cond_33_shl = {mux_cond_33, 1'h0};
  assign mux_cond_33_pad = {18'h0,mux_cond_33_shl};
  assign mux_cond_34_shl = {mux_cond_34, 1'h0};
  assign mux_cond_34_pad = {18'h0,mux_cond_34_shl};
  assign mux_cond_35_shl = {mux_cond_35, 3'h0};
  assign mux_cond_35_pad = {16'h0,mux_cond_35_shl};
  assign mux_cond_36_shl = {mux_cond_36, 7'h0};
  assign mux_cond_36_pad = {12'h0,mux_cond_36_shl};
  assign mux_cond_37_shl = {mux_cond_37, 6'h0};
  assign mux_cond_37_pad = {13'h0,mux_cond_37_shl};
  assign mux_cond_38_shl = {mux_cond_38, 5'h0};
  assign mux_cond_38_pad = {14'h0,mux_cond_38_shl};
  assign mux_cond_39_shl = {mux_cond_39, 4'h0};
  assign mux_cond_39_pad = {15'h0,mux_cond_39_shl};
  assign mux_cond_40_shl = {mux_cond_40, 3'h0};
  assign mux_cond_40_pad = {16'h0,mux_cond_40_shl};
  assign mux_cond_41_shl = {mux_cond_41, 10'h0};
  assign mux_cond_41_pad = {9'h0,mux_cond_41_shl};
  assign mux_cond_42_shl = {mux_cond_42, 14'h0};
  assign mux_cond_42_pad = {5'h0,mux_cond_42_shl};
  assign mux_cond_43_shl = {mux_cond_43, 16'h0};
  assign mux_cond_43_pad = {3'h0,mux_cond_43_shl};
  assign mux_cond_44_shl = {mux_cond_44, 2'h0};
  assign mux_cond_44_pad = {17'h0,mux_cond_44_shl};
  assign mux_cond_45_shl = {mux_cond_45, 13'h0};
  assign mux_cond_45_pad = {6'h0,mux_cond_45_shl};
  assign mux_cond_46_shl = {mux_cond_46, 4'h0};
  assign mux_cond_46_pad = {15'h0,mux_cond_46_shl};
  assign mux_cond_47_shl = {mux_cond_47, 8'h0};
  assign mux_cond_47_pad = {11'h0,mux_cond_47_shl};
  assign mux_cond_48_shl = {mux_cond_48, 10'h0};
  assign mux_cond_48_pad = {9'h0,mux_cond_48_shl};
  assign mux_cond_49_shl = {mux_cond_49, 8'h0};
  assign mux_cond_49_pad = {11'h0,mux_cond_49_shl};
  assign mux_cond_50_shl = {mux_cond_50, 16'h0};
  assign mux_cond_50_pad = {3'h0,mux_cond_50_shl};
  assign mux_cond_51_shl = {mux_cond_51, 12'h0};
  assign mux_cond_51_pad = {7'h0,mux_cond_51_shl};
  assign mux_cond_52_shl = {mux_cond_52, 19'h0};
  assign mux_cond_52_pad = mux_cond_52_shl;
  assign mux_cond_53_shl = {mux_cond_53, 16'h0};
  assign mux_cond_53_pad = {3'h0,mux_cond_53_shl};
  assign mux_cond_54_shl = {mux_cond_54, 19'h0};
  assign mux_cond_54_pad = mux_cond_54_shl;
  assign mux_cond_55_shl = {mux_cond_55, 10'h0};
  assign mux_cond_55_pad = {9'h0,mux_cond_55_shl};
  assign mux_cond_56_shl = {mux_cond_56, 7'h0};
  assign mux_cond_56_pad = {12'h0,mux_cond_56_shl};
  assign mux_cond_57_shl = {mux_cond_57, 1'h0};
  assign mux_cond_57_pad = {18'h0,mux_cond_57_shl};
  assign mux_cond_58_shl = {mux_cond_58, 13'h0};
  assign mux_cond_58_pad = {6'h0,mux_cond_58_shl};
  assign mux_cond_59_shl = {mux_cond_59, 18'h0};
  assign mux_cond_59_pad = {1'h0,mux_cond_59_shl};
  assign mux_cond_60_shl = {mux_cond_60, 14'h0};
  assign mux_cond_60_pad = {5'h0,mux_cond_60_shl};
  assign mux_cond_61_shl = {mux_cond_61, 2'h0};
  assign mux_cond_61_pad = {17'h0,mux_cond_61_shl};
  assign mux_cond_62_shl = {mux_cond_62, 17'h0};
  assign mux_cond_62_pad = {2'h0,mux_cond_62_shl};
  assign mux_cond_63_shl = {mux_cond_63, 3'h0};
  assign mux_cond_63_pad = {16'h0,mux_cond_63_shl};
  assign mux_cond_64_shl = {mux_cond_64, 14'h0};
  assign mux_cond_64_pad = {5'h0,mux_cond_64_shl};
  assign mux_cond_65_shl = {mux_cond_65, 7'h0};
  assign mux_cond_65_pad = {12'h0,mux_cond_65_shl};
  assign mux_cond_66_shl = {mux_cond_66, 15'h0};
  assign mux_cond_66_pad = {4'h0,mux_cond_66_shl};
  assign mux_cond_67_shl = {mux_cond_67, 16'h0};
  assign mux_cond_67_pad = {3'h0,mux_cond_67_shl};
  assign mux_cond_68_shl = {mux_cond_68, 12'h0};
  assign mux_cond_68_pad = {7'h0,mux_cond_68_shl};
  assign mux_cond_69_shl = {mux_cond_69, 1'h0};
  assign mux_cond_69_pad = {18'h0,mux_cond_69_shl};
  assign mux_cond_70_shl = {mux_cond_70, 5'h0};
  assign mux_cond_70_pad = {14'h0,mux_cond_70_shl};
  assign mux_cond_71_shl = {mux_cond_71, 11'h0};
  assign mux_cond_71_pad = {8'h0,mux_cond_71_shl};
  assign mux_cond_72_shl = {mux_cond_72, 13'h0};
  assign mux_cond_72_pad = {6'h0,mux_cond_72_shl};
  assign mux_cond_73_shl = {mux_cond_73, 13'h0};
  assign mux_cond_73_pad = {6'h0,mux_cond_73_shl};
  assign sectored_entries_7_valid_1_shl = {sectored_entries_7_valid_1, 2'h0};
  assign sectored_entries_7_valid_1_pad = {17'h0,sectored_entries_7_valid_1_shl};
  assign sectored_entries_5_valid_3_shl = {sectored_entries_5_valid_3, 13'h0};
  assign sectored_entries_5_valid_3_pad = {6'h0,sectored_entries_5_valid_3_shl};
  assign sectored_entries_5_valid_1_shl = {sectored_entries_5_valid_1, 2'h0};
  assign sectored_entries_5_valid_1_pad = {17'h0,sectored_entries_5_valid_1_shl};
  assign sectored_entries_4_valid_1_shl = {sectored_entries_4_valid_1, 2'h0};
  assign sectored_entries_4_valid_1_pad = {17'h0,sectored_entries_4_valid_1_shl};
  assign superpage_entries_0_valid_0_shl = {superpage_entries_0_valid_0, 5'h0};
  assign superpage_entries_0_valid_0_pad = {14'h0,superpage_entries_0_valid_0_shl};
  assign sectored_entries_3_valid_2_shl = {sectored_entries_3_valid_2, 17'h0};
  assign sectored_entries_3_valid_2_pad = {2'h0,sectored_entries_3_valid_2_shl};
  assign sectored_entries_1_valid_0_shl = {sectored_entries_1_valid_0, 17'h0};
  assign sectored_entries_1_valid_0_pad = {2'h0,sectored_entries_1_valid_0_shl};
  assign superpage_entries_3_level_shl = {superpage_entries_3_level, 10'h0};
  assign superpage_entries_3_level_pad = {8'h0,superpage_entries_3_level_shl};
  assign sectored_entries_5_valid_0_shl = {sectored_entries_5_valid_0, 17'h0};
  assign sectored_entries_5_valid_0_pad = {2'h0,sectored_entries_5_valid_0_shl};
  assign sectored_entries_0_valid_1_shl = {sectored_entries_0_valid_1, 2'h0};
  assign sectored_entries_0_valid_1_pad = {17'h0,sectored_entries_0_valid_1_shl};
  assign sectored_entries_3_valid_0_shl = {sectored_entries_3_valid_0, 17'h0};
  assign sectored_entries_3_valid_0_pad = {2'h0,sectored_entries_3_valid_0_shl};
  assign sectored_entries_7_valid_2_shl = {sectored_entries_7_valid_2, 17'h0};
  assign sectored_entries_7_valid_2_pad = {2'h0,sectored_entries_7_valid_2_shl};
  assign sectored_entries_2_valid_3_shl = {sectored_entries_2_valid_3, 13'h0};
  assign sectored_entries_2_valid_3_pad = {6'h0,sectored_entries_2_valid_3_shl};
  assign sectored_entries_4_valid_0_shl = {sectored_entries_4_valid_0, 17'h0};
  assign sectored_entries_4_valid_0_pad = {2'h0,sectored_entries_4_valid_0_shl};
  assign sectored_entries_6_valid_3_shl = {sectored_entries_6_valid_3, 13'h0};
  assign sectored_entries_6_valid_3_pad = {6'h0,sectored_entries_6_valid_3_shl};
  assign sectored_entries_1_valid_3_shl = {sectored_entries_1_valid_3, 13'h0};
  assign sectored_entries_1_valid_3_pad = {6'h0,sectored_entries_1_valid_3_shl};
  assign sectored_entries_6_valid_0_shl = {sectored_entries_6_valid_0, 17'h0};
  assign sectored_entries_6_valid_0_pad = {2'h0,sectored_entries_6_valid_0_shl};
  assign sectored_entries_2_valid_2_shl = {sectored_entries_2_valid_2, 17'h0};
  assign sectored_entries_2_valid_2_pad = {2'h0,sectored_entries_2_valid_2_shl};
  assign sectored_entries_6_valid_2_shl = {sectored_entries_6_valid_2, 17'h0};
  assign sectored_entries_6_valid_2_pad = {2'h0,sectored_entries_6_valid_2_shl};
  assign sectored_entries_6_valid_1_shl = {sectored_entries_6_valid_1, 2'h0};
  assign sectored_entries_6_valid_1_pad = {17'h0,sectored_entries_6_valid_1_shl};
  assign sectored_entries_4_valid_3_shl = {sectored_entries_4_valid_3, 13'h0};
  assign sectored_entries_4_valid_3_pad = {6'h0,sectored_entries_4_valid_3_shl};
  assign sectored_entries_1_valid_2_shl = {sectored_entries_1_valid_2, 17'h0};
  assign sectored_entries_1_valid_2_pad = {2'h0,sectored_entries_1_valid_2_shl};
  assign sectored_entries_5_valid_2_shl = {sectored_entries_5_valid_2, 17'h0};
  assign sectored_entries_5_valid_2_pad = {2'h0,sectored_entries_5_valid_2_shl};
  assign superpage_entries_2_level_shl = {superpage_entries_2_level, 10'h0};
  assign superpage_entries_2_level_pad = {8'h0,superpage_entries_2_level_shl};
  assign superpage_entries_3_valid_0_shl = {superpage_entries_3_valid_0, 5'h0};
  assign superpage_entries_3_valid_0_pad = {14'h0,superpage_entries_3_valid_0_shl};
  assign sectored_entries_1_valid_1_shl = {sectored_entries_1_valid_1, 2'h0};
  assign sectored_entries_1_valid_1_pad = {17'h0,sectored_entries_1_valid_1_shl};
  assign sectored_entries_0_valid_0_shl = {sectored_entries_0_valid_0, 17'h0};
  assign sectored_entries_0_valid_0_pad = {2'h0,sectored_entries_0_valid_0_shl};
  assign superpage_entries_1_valid_0_shl = {superpage_entries_1_valid_0, 5'h0};
  assign superpage_entries_1_valid_0_pad = {14'h0,superpage_entries_1_valid_0_shl};
  assign sectored_entries_0_valid_3_shl = {sectored_entries_0_valid_3, 13'h0};
  assign sectored_entries_0_valid_3_pad = {6'h0,sectored_entries_0_valid_3_shl};
  assign sectored_entries_7_valid_0_shl = {sectored_entries_7_valid_0, 17'h0};
  assign sectored_entries_7_valid_0_pad = {2'h0,sectored_entries_7_valid_0_shl};
  assign sectored_entries_0_valid_2_shl = {sectored_entries_0_valid_2, 17'h0};
  assign sectored_entries_0_valid_2_pad = {2'h0,sectored_entries_0_valid_2_shl};
  assign superpage_entries_0_level_shl = {superpage_entries_0_level, 10'h0};
  assign superpage_entries_0_level_pad = {8'h0,superpage_entries_0_level_shl};
  assign sectored_entries_2_valid_1_shl = {sectored_entries_2_valid_1, 2'h0};
  assign sectored_entries_2_valid_1_pad = {17'h0,sectored_entries_2_valid_1_shl};
  assign sectored_entries_3_valid_1_shl = {sectored_entries_3_valid_1, 2'h0};
  assign sectored_entries_3_valid_1_pad = {17'h0,sectored_entries_3_valid_1_shl};
  assign sectored_entries_2_valid_0_shl = {sectored_entries_2_valid_0, 17'h0};
  assign sectored_entries_2_valid_0_pad = {2'h0,sectored_entries_2_valid_0_shl};
  assign sectored_entries_7_valid_3_shl = {sectored_entries_7_valid_3, 13'h0};
  assign sectored_entries_7_valid_3_pad = {6'h0,sectored_entries_7_valid_3_shl};
  assign sectored_entries_4_valid_2_shl = {sectored_entries_4_valid_2, 17'h0};
  assign sectored_entries_4_valid_2_pad = {2'h0,sectored_entries_4_valid_2_shl};
  assign sectored_entries_3_valid_3_shl = {sectored_entries_3_valid_3, 13'h0};
  assign sectored_entries_3_valid_3_pad = {6'h0,sectored_entries_3_valid_3_shl};
  assign superpage_entries_1_level_shl = {superpage_entries_1_level, 10'h0};
  assign superpage_entries_1_level_pad = {8'h0,superpage_entries_1_level_shl};
  assign superpage_entries_2_valid_0_shl = {superpage_entries_2_valid_0, 5'h0};
  assign superpage_entries_2_valid_0_pad = {14'h0,superpage_entries_2_valid_0_shl};
  assign TLB_xor64 = state_pad ^ r_sectored_repl_addr_pad;
  assign TLB_xor31 = r_superpage_repl_addr_pad ^ TLB_xor64;
  assign TLB_xor65 = r_sectored_hit_addr_pad ^ special_entry_valid_0_pad;
  assign TLB_xor66 = special_entry_level_pad ^ r_sectored_hit_pad;
  assign TLB_xor32 = TLB_xor65 ^ TLB_xor66;
  assign TLB_xor15 = TLB_xor31 ^ TLB_xor32;
  assign TLB_xor67 = mux_cond_0_pad ^ mux_cond_1_pad;
  assign TLB_xor68 = mux_cond_2_pad ^ mux_cond_3_pad;
  assign TLB_xor33 = TLB_xor67 ^ TLB_xor68;
  assign TLB_xor69 = mux_cond_4_pad ^ mux_cond_5_pad;
  assign TLB_xor70 = mux_cond_6_pad ^ mux_cond_7_pad;
  assign TLB_xor34 = TLB_xor69 ^ TLB_xor70;
  assign TLB_xor16 = TLB_xor33 ^ TLB_xor34;
  assign TLB_xor7 = TLB_xor15 ^ TLB_xor16;
  assign TLB_xor72 = mux_cond_9_pad ^ mux_cond_10_pad;
  assign TLB_xor35 = mux_cond_8_pad ^ TLB_xor72;
  assign TLB_xor73 = mux_cond_11_pad ^ mux_cond_12_pad;
  assign TLB_xor74 = mux_cond_13_pad ^ mux_cond_14_pad;
  assign TLB_xor36 = TLB_xor73 ^ TLB_xor74;
  assign TLB_xor17 = TLB_xor35 ^ TLB_xor36;
  assign TLB_xor75 = mux_cond_15_pad ^ mux_cond_16_pad;
  assign TLB_xor76 = mux_cond_17_pad ^ mux_cond_18_pad;
  assign TLB_xor37 = TLB_xor75 ^ TLB_xor76;
  assign TLB_xor77 = mux_cond_19_pad ^ mux_cond_20_pad;
  assign TLB_xor78 = mux_cond_21_pad ^ mux_cond_22_pad;
  assign TLB_xor38 = TLB_xor77 ^ TLB_xor78;
  assign TLB_xor18 = TLB_xor37 ^ TLB_xor38;
  assign TLB_xor8 = TLB_xor17 ^ TLB_xor18;
  assign TLB_xor3 = TLB_xor7 ^ TLB_xor8;
  assign TLB_xor80 = mux_cond_24_pad ^ mux_cond_25_pad;
  assign TLB_xor39 = mux_cond_23_pad ^ TLB_xor80;
  assign TLB_xor81 = mux_cond_26_pad ^ mux_cond_27_pad;
  assign TLB_xor82 = mux_cond_28_pad ^ mux_cond_29_pad;
  assign TLB_xor40 = TLB_xor81 ^ TLB_xor82;
  assign TLB_xor19 = TLB_xor39 ^ TLB_xor40;
  assign TLB_xor83 = mux_cond_30_pad ^ mux_cond_31_pad;
  assign TLB_xor84 = mux_cond_32_pad ^ mux_cond_33_pad;
  assign TLB_xor41 = TLB_xor83 ^ TLB_xor84;
  assign TLB_xor85 = mux_cond_34_pad ^ mux_cond_35_pad;
  assign TLB_xor86 = mux_cond_36_pad ^ mux_cond_37_pad;
  assign TLB_xor42 = TLB_xor85 ^ TLB_xor86;
  assign TLB_xor20 = TLB_xor41 ^ TLB_xor42;
  assign TLB_xor9 = TLB_xor19 ^ TLB_xor20;
  assign TLB_xor88 = mux_cond_39_pad ^ mux_cond_40_pad;
  assign TLB_xor43 = mux_cond_38_pad ^ TLB_xor88;
  assign TLB_xor89 = mux_cond_41_pad ^ mux_cond_42_pad;
  assign TLB_xor90 = mux_cond_43_pad ^ mux_cond_44_pad;
  assign TLB_xor44 = TLB_xor89 ^ TLB_xor90;
  assign TLB_xor21 = TLB_xor43 ^ TLB_xor44;
  assign TLB_xor91 = mux_cond_45_pad ^ mux_cond_46_pad;
  assign TLB_xor92 = mux_cond_47_pad ^ mux_cond_48_pad;
  assign TLB_xor45 = TLB_xor91 ^ TLB_xor92;
  assign TLB_xor93 = mux_cond_49_pad ^ mux_cond_50_pad;
  assign TLB_xor94 = mux_cond_51_pad ^ mux_cond_52_pad;
  assign TLB_xor46 = TLB_xor93 ^ TLB_xor94;
  assign TLB_xor22 = TLB_xor45 ^ TLB_xor46;
  assign TLB_xor10 = TLB_xor21 ^ TLB_xor22;
  assign TLB_xor4 = TLB_xor9 ^ TLB_xor10;
  assign TLB_xor1 = TLB_xor3 ^ TLB_xor4;
  assign TLB_xor96 = mux_cond_54_pad ^ mux_cond_55_pad;
  assign TLB_xor47 = mux_cond_53_pad ^ TLB_xor96;
  assign TLB_xor97 = mux_cond_56_pad ^ mux_cond_57_pad;
  assign TLB_xor98 = mux_cond_58_pad ^ mux_cond_59_pad;
  assign TLB_xor48 = TLB_xor97 ^ TLB_xor98;
  assign TLB_xor23 = TLB_xor47 ^ TLB_xor48;
  assign TLB_xor99 = mux_cond_60_pad ^ mux_cond_61_pad;
  assign TLB_xor100 = mux_cond_62_pad ^ mux_cond_63_pad;
  assign TLB_xor49 = TLB_xor99 ^ TLB_xor100;
  assign TLB_xor101 = mux_cond_64_pad ^ mux_cond_65_pad;
  assign TLB_xor102 = mux_cond_66_pad ^ mux_cond_67_pad;
  assign TLB_xor50 = TLB_xor101 ^ TLB_xor102;
  assign TLB_xor24 = TLB_xor49 ^ TLB_xor50;
  assign TLB_xor11 = TLB_xor23 ^ TLB_xor24;
  assign TLB_xor104 = mux_cond_69_pad ^ mux_cond_70_pad;
  assign TLB_xor51 = mux_cond_68_pad ^ TLB_xor104;
  assign TLB_xor105 = mux_cond_71_pad ^ mux_cond_72_pad;
  assign TLB_xor106 = mux_cond_73_pad ^ sectored_entries_7_valid_1_pad;
  assign TLB_xor52 = TLB_xor105 ^ TLB_xor106;
  assign TLB_xor25 = TLB_xor51 ^ TLB_xor52;
  assign TLB_xor107 = sectored_entries_5_valid_3_pad ^ sectored_entries_5_valid_1_pad;
  assign TLB_xor108 = sectored_entries_4_valid_1_pad ^ superpage_entries_0_valid_0_pad;
  assign TLB_xor53 = TLB_xor107 ^ TLB_xor108;
  assign TLB_xor109 = sectored_entries_3_valid_2_pad ^ sectored_entries_1_valid_0_pad;
  assign TLB_xor110 = superpage_entries_3_level_pad ^ sectored_entries_5_valid_0_pad;
  assign TLB_xor54 = TLB_xor109 ^ TLB_xor110;
  assign TLB_xor26 = TLB_xor53 ^ TLB_xor54;
  assign TLB_xor12 = TLB_xor25 ^ TLB_xor26;
  assign TLB_xor5 = TLB_xor11 ^ TLB_xor12;
  assign TLB_xor112 = sectored_entries_3_valid_0_pad ^ sectored_entries_7_valid_2_pad;
  assign TLB_xor55 = sectored_entries_0_valid_1_pad ^ TLB_xor112;
  assign TLB_xor113 = sectored_entries_2_valid_3_pad ^ sectored_entries_4_valid_0_pad;
  assign TLB_xor114 = sectored_entries_6_valid_3_pad ^ sectored_entries_1_valid_3_pad;
  assign TLB_xor56 = TLB_xor113 ^ TLB_xor114;
  assign TLB_xor27 = TLB_xor55 ^ TLB_xor56;
  assign TLB_xor115 = sectored_entries_6_valid_0_pad ^ sectored_entries_2_valid_2_pad;
  assign TLB_xor116 = sectored_entries_6_valid_2_pad ^ sectored_entries_6_valid_1_pad;
  assign TLB_xor57 = TLB_xor115 ^ TLB_xor116;
  assign TLB_xor117 = sectored_entries_4_valid_3_pad ^ sectored_entries_1_valid_2_pad;
  assign TLB_xor118 = sectored_entries_5_valid_2_pad ^ superpage_entries_2_level_pad;
  assign TLB_xor58 = TLB_xor117 ^ TLB_xor118;
  assign TLB_xor28 = TLB_xor57 ^ TLB_xor58;
  assign TLB_xor13 = TLB_xor27 ^ TLB_xor28;
  assign TLB_xor119 = superpage_entries_3_valid_0_pad ^ sectored_entries_1_valid_1_pad;
  assign TLB_xor120 = sectored_entries_0_valid_0_pad ^ superpage_entries_1_valid_0_pad;
  assign TLB_xor59 = TLB_xor119 ^ TLB_xor120;
  assign TLB_xor121 = sectored_entries_0_valid_3_pad ^ sectored_entries_7_valid_0_pad;
  assign TLB_xor122 = sectored_entries_0_valid_2_pad ^ superpage_entries_0_level_pad;
  assign TLB_xor60 = TLB_xor121 ^ TLB_xor122;
  assign TLB_xor29 = TLB_xor59 ^ TLB_xor60;
  assign TLB_xor123 = sectored_entries_2_valid_1_pad ^ sectored_entries_3_valid_1_pad;
  assign TLB_xor124 = sectored_entries_2_valid_0_pad ^ sectored_entries_7_valid_3_pad;
  assign TLB_xor61 = TLB_xor123 ^ TLB_xor124;
  assign TLB_xor125 = sectored_entries_4_valid_2_pad ^ sectored_entries_3_valid_3_pad;
  assign TLB_xor126 = superpage_entries_1_level_pad ^ superpage_entries_2_valid_0_pad;
  assign TLB_xor62 = TLB_xor125 ^ TLB_xor126;
  assign TLB_xor30 = TLB_xor61 ^ TLB_xor62;
  assign TLB_xor14 = TLB_xor29 ^ TLB_xor30;
  assign TLB_xor6 = TLB_xor13 ^ TLB_xor14;
  assign TLB_xor2 = TLB_xor5 ^ TLB_xor6;
  assign TLB_xor0 = TLB_xor1 ^ TLB_xor2;
  assign pmp_sum = TLB_covSum + pmp_io_covSum;
  assign io_covSum = pmp_sum;
  assign stopEn0 = io_sfence_valid & ~_T_2949;
  assign pmp_metaAssert_wire = pmp_metaAssert;
  assign TLB_or0 = stopEn0 | pmp_metaAssert_wire;
  assign metaAssert = TLB_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sectored_entries_0_tag = _RAND_0[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  sectored_entries_0_data_0 = _RAND_1[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  sectored_entries_0_data_1 = _RAND_2[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{`RANDOM}};
  sectored_entries_0_data_2 = _RAND_3[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{`RANDOM}};
  sectored_entries_0_data_3 = _RAND_4[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  sectored_entries_0_valid_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sectored_entries_0_valid_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  sectored_entries_0_valid_2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sectored_entries_0_valid_3 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  sectored_entries_1_tag = _RAND_9[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {2{`RANDOM}};
  sectored_entries_1_data_0 = _RAND_10[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{`RANDOM}};
  sectored_entries_1_data_1 = _RAND_11[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {2{`RANDOM}};
  sectored_entries_1_data_2 = _RAND_12[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  sectored_entries_1_data_3 = _RAND_13[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  sectored_entries_1_valid_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  sectored_entries_1_valid_1 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  sectored_entries_1_valid_2 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  sectored_entries_1_valid_3 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  sectored_entries_2_tag = _RAND_18[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{`RANDOM}};
  sectored_entries_2_data_0 = _RAND_19[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{`RANDOM}};
  sectored_entries_2_data_1 = _RAND_20[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{`RANDOM}};
  sectored_entries_2_data_2 = _RAND_21[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {2{`RANDOM}};
  sectored_entries_2_data_3 = _RAND_22[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  sectored_entries_2_valid_0 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  sectored_entries_2_valid_1 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  sectored_entries_2_valid_2 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  sectored_entries_2_valid_3 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  sectored_entries_3_tag = _RAND_27[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {2{`RANDOM}};
  sectored_entries_3_data_0 = _RAND_28[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {2{`RANDOM}};
  sectored_entries_3_data_1 = _RAND_29[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {2{`RANDOM}};
  sectored_entries_3_data_2 = _RAND_30[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{`RANDOM}};
  sectored_entries_3_data_3 = _RAND_31[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  sectored_entries_3_valid_0 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  sectored_entries_3_valid_1 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  sectored_entries_3_valid_2 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  sectored_entries_3_valid_3 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  sectored_entries_4_tag = _RAND_36[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{`RANDOM}};
  sectored_entries_4_data_0 = _RAND_37[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {2{`RANDOM}};
  sectored_entries_4_data_1 = _RAND_38[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{`RANDOM}};
  sectored_entries_4_data_2 = _RAND_39[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {2{`RANDOM}};
  sectored_entries_4_data_3 = _RAND_40[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  sectored_entries_4_valid_0 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  sectored_entries_4_valid_1 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  sectored_entries_4_valid_2 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  sectored_entries_4_valid_3 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  sectored_entries_5_tag = _RAND_45[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {2{`RANDOM}};
  sectored_entries_5_data_0 = _RAND_46[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {2{`RANDOM}};
  sectored_entries_5_data_1 = _RAND_47[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {2{`RANDOM}};
  sectored_entries_5_data_2 = _RAND_48[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {2{`RANDOM}};
  sectored_entries_5_data_3 = _RAND_49[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  sectored_entries_5_valid_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  sectored_entries_5_valid_1 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  sectored_entries_5_valid_2 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  sectored_entries_5_valid_3 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  sectored_entries_6_tag = _RAND_54[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {2{`RANDOM}};
  sectored_entries_6_data_0 = _RAND_55[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {2{`RANDOM}};
  sectored_entries_6_data_1 = _RAND_56[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {2{`RANDOM}};
  sectored_entries_6_data_2 = _RAND_57[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {2{`RANDOM}};
  sectored_entries_6_data_3 = _RAND_58[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  sectored_entries_6_valid_0 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  sectored_entries_6_valid_1 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  sectored_entries_6_valid_2 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  sectored_entries_6_valid_3 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  sectored_entries_7_tag = _RAND_63[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {2{`RANDOM}};
  sectored_entries_7_data_0 = _RAND_64[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {2{`RANDOM}};
  sectored_entries_7_data_1 = _RAND_65[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {2{`RANDOM}};
  sectored_entries_7_data_2 = _RAND_66[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {2{`RANDOM}};
  sectored_entries_7_data_3 = _RAND_67[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  sectored_entries_7_valid_0 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  sectored_entries_7_valid_1 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  sectored_entries_7_valid_2 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  sectored_entries_7_valid_3 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  superpage_entries_0_level = _RAND_72[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  superpage_entries_0_tag = _RAND_73[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {2{`RANDOM}};
  superpage_entries_0_data_0 = _RAND_74[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  superpage_entries_0_valid_0 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  superpage_entries_1_level = _RAND_76[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  superpage_entries_1_tag = _RAND_77[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {2{`RANDOM}};
  superpage_entries_1_data_0 = _RAND_78[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  superpage_entries_1_valid_0 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  superpage_entries_2_level = _RAND_80[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  superpage_entries_2_tag = _RAND_81[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {2{`RANDOM}};
  superpage_entries_2_data_0 = _RAND_82[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  superpage_entries_2_valid_0 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  superpage_entries_3_level = _RAND_84[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  superpage_entries_3_tag = _RAND_85[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {2{`RANDOM}};
  superpage_entries_3_data_0 = _RAND_86[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  superpage_entries_3_valid_0 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  special_entry_level = _RAND_88[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  special_entry_tag = _RAND_89[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {2{`RANDOM}};
  special_entry_data_0 = _RAND_90[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  special_entry_valid_0 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  state = _RAND_92[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  r_refill_tag = _RAND_93[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  r_superpage_repl_addr = _RAND_94[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  r_sectored_repl_addr = _RAND_95[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  r_sectored_hit_addr = _RAND_96[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  r_sectored_hit = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  vpoffset_cfg_value = _RAND_98[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  requestedVPN = _RAND_99[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_2554 = _RAND_100[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_2556 = _RAND_101[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  TLB_state = _RAND_102[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    TLB_cov[initvar] = _RAND_103[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  TLB_covSum = _RAND_104[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  TLB_metaAssert = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      sectored_entries_0_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1505) begin
            sectored_entries_0_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1505) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_0 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_data_1 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1505) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_1 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_data_2 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1505) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_2 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_data_3 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1505) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_3 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_0_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2957) begin
          if (sectored_entries_0_data_0[0]) begin
            sectored_entries_0_valid_0 <= 1'h0;
          end else if (_T_727) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_0_valid_0 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1505) begin
                    sectored_entries_0_valid_0 <= _GEN_85;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1505) begin
                  sectored_entries_0_valid_0 <= _GEN_85;
                end
              end
            end
          end
        end else if (_T_727) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_0_valid_0 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1505) begin
                  sectored_entries_0_valid_0 <= _GEN_85;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1505) begin
                sectored_entries_0_valid_0 <= _GEN_85;
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_0 <= _GEN_656;
      end
    end else begin
      sectored_entries_0_valid_0 <= _GEN_473;
    end
    if (metaReset) begin
      sectored_entries_0_valid_1 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_0_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2957) begin
          if (sectored_entries_0_data_1[0]) begin
            sectored_entries_0_valid_1 <= 1'h0;
          end else if (_T_727) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_0_valid_1 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1505) begin
                    sectored_entries_0_valid_1 <= _GEN_86;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1505) begin
                  sectored_entries_0_valid_1 <= _GEN_86;
                end
              end
            end
          end
        end else if (_T_727) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_0_valid_1 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1505) begin
                  sectored_entries_0_valid_1 <= _GEN_86;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1505) begin
                sectored_entries_0_valid_1 <= _GEN_86;
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_1 <= _GEN_657;
      end
    end else begin
      sectored_entries_0_valid_1 <= _GEN_474;
    end
    if (metaReset) begin
      sectored_entries_0_valid_2 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_0_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2957) begin
          if (sectored_entries_0_data_2[0]) begin
            sectored_entries_0_valid_2 <= 1'h0;
          end else if (_T_727) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_0_valid_2 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1505) begin
                    sectored_entries_0_valid_2 <= _GEN_87;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1505) begin
                  sectored_entries_0_valid_2 <= _GEN_87;
                end
              end
            end
          end
        end else if (_T_727) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_0_valid_2 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1505) begin
                  sectored_entries_0_valid_2 <= _GEN_87;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1505) begin
                sectored_entries_0_valid_2 <= _GEN_87;
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_2 <= _GEN_658;
      end
    end else begin
      sectored_entries_0_valid_2 <= _GEN_475;
    end
    if (metaReset) begin
      sectored_entries_0_valid_3 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_0_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2957) begin
          if (sectored_entries_0_data_3[0]) begin
            sectored_entries_0_valid_3 <= 1'h0;
          end else if (_T_727) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_0_valid_3 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1505) begin
                    sectored_entries_0_valid_3 <= _GEN_88;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1505) begin
                  sectored_entries_0_valid_3 <= _GEN_88;
                end
              end
            end
          end
        end else if (_T_727) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_0_valid_3 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1505) begin
                  sectored_entries_0_valid_3 <= _GEN_88;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1505) begin
                sectored_entries_0_valid_3 <= _GEN_88;
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_3 <= _GEN_659;
      end
    end else begin
      sectored_entries_0_valid_3 <= _GEN_476;
    end
    if (metaReset) begin
      sectored_entries_1_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1522) begin
            sectored_entries_1_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_1_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1522) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_0 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_1_data_1 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1522) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_1 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_1_data_2 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1522) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_2 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_1_data_3 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1522) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_3 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_1_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_1_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3128) begin
          if (sectored_entries_1_data_0[0]) begin
            sectored_entries_1_valid_0 <= 1'h0;
          end else if (_T_733) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_1_valid_0 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1522) begin
                    sectored_entries_1_valid_0 <= _GEN_107;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1522) begin
                  sectored_entries_1_valid_0 <= _GEN_107;
                end
              end
            end
          end
        end else if (_T_733) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_1_valid_0 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1522) begin
                  sectored_entries_1_valid_0 <= _GEN_107;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1522) begin
                sectored_entries_1_valid_0 <= _GEN_107;
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_0 <= _GEN_684;
      end
    end else begin
      sectored_entries_1_valid_0 <= _GEN_483;
    end
    if (metaReset) begin
      sectored_entries_1_valid_1 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_1_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3128) begin
          if (sectored_entries_1_data_1[0]) begin
            sectored_entries_1_valid_1 <= 1'h0;
          end else if (_T_733) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_1_valid_1 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1522) begin
                    sectored_entries_1_valid_1 <= _GEN_108;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1522) begin
                  sectored_entries_1_valid_1 <= _GEN_108;
                end
              end
            end
          end
        end else if (_T_733) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_1_valid_1 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1522) begin
                  sectored_entries_1_valid_1 <= _GEN_108;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1522) begin
                sectored_entries_1_valid_1 <= _GEN_108;
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_1 <= _GEN_685;
      end
    end else begin
      sectored_entries_1_valid_1 <= _GEN_484;
    end
    if (metaReset) begin
      sectored_entries_1_valid_2 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_1_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3128) begin
          if (sectored_entries_1_data_2[0]) begin
            sectored_entries_1_valid_2 <= 1'h0;
          end else if (_T_733) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_1_valid_2 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1522) begin
                    sectored_entries_1_valid_2 <= _GEN_109;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1522) begin
                  sectored_entries_1_valid_2 <= _GEN_109;
                end
              end
            end
          end
        end else if (_T_733) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_1_valid_2 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1522) begin
                  sectored_entries_1_valid_2 <= _GEN_109;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1522) begin
                sectored_entries_1_valid_2 <= _GEN_109;
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_2 <= _GEN_686;
      end
    end else begin
      sectored_entries_1_valid_2 <= _GEN_485;
    end
    if (metaReset) begin
      sectored_entries_1_valid_3 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_1_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3128) begin
          if (sectored_entries_1_data_3[0]) begin
            sectored_entries_1_valid_3 <= 1'h0;
          end else if (_T_733) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_1_valid_3 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1522) begin
                    sectored_entries_1_valid_3 <= _GEN_110;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1522) begin
                  sectored_entries_1_valid_3 <= _GEN_110;
                end
              end
            end
          end
        end else if (_T_733) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_1_valid_3 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1522) begin
                  sectored_entries_1_valid_3 <= _GEN_110;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1522) begin
                sectored_entries_1_valid_3 <= _GEN_110;
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_3 <= _GEN_687;
      end
    end else begin
      sectored_entries_1_valid_3 <= _GEN_486;
    end
    if (metaReset) begin
      sectored_entries_2_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1539) begin
            sectored_entries_2_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_2_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1539) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_0 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_2_data_1 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1539) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_1 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_2_data_2 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1539) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_2 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_2_data_3 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1539) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_3 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_2_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_2_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3299) begin
          if (sectored_entries_2_data_0[0]) begin
            sectored_entries_2_valid_0 <= 1'h0;
          end else if (_T_739) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_2_valid_0 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1539) begin
                    sectored_entries_2_valid_0 <= _GEN_129;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1539) begin
                  sectored_entries_2_valid_0 <= _GEN_129;
                end
              end
            end
          end
        end else if (_T_739) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_2_valid_0 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1539) begin
                  sectored_entries_2_valid_0 <= _GEN_129;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1539) begin
                sectored_entries_2_valid_0 <= _GEN_129;
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_0 <= _GEN_712;
      end
    end else begin
      sectored_entries_2_valid_0 <= _GEN_493;
    end
    if (metaReset) begin
      sectored_entries_2_valid_1 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_2_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3299) begin
          if (sectored_entries_2_data_1[0]) begin
            sectored_entries_2_valid_1 <= 1'h0;
          end else if (_T_739) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_2_valid_1 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1539) begin
                    sectored_entries_2_valid_1 <= _GEN_130;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1539) begin
                  sectored_entries_2_valid_1 <= _GEN_130;
                end
              end
            end
          end
        end else if (_T_739) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_2_valid_1 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1539) begin
                  sectored_entries_2_valid_1 <= _GEN_130;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1539) begin
                sectored_entries_2_valid_1 <= _GEN_130;
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_1 <= _GEN_713;
      end
    end else begin
      sectored_entries_2_valid_1 <= _GEN_494;
    end
    if (metaReset) begin
      sectored_entries_2_valid_2 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_2_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3299) begin
          if (sectored_entries_2_data_2[0]) begin
            sectored_entries_2_valid_2 <= 1'h0;
          end else if (_T_739) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_2_valid_2 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1539) begin
                    sectored_entries_2_valid_2 <= _GEN_131;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1539) begin
                  sectored_entries_2_valid_2 <= _GEN_131;
                end
              end
            end
          end
        end else if (_T_739) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_2_valid_2 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1539) begin
                  sectored_entries_2_valid_2 <= _GEN_131;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1539) begin
                sectored_entries_2_valid_2 <= _GEN_131;
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_2 <= _GEN_714;
      end
    end else begin
      sectored_entries_2_valid_2 <= _GEN_495;
    end
    if (metaReset) begin
      sectored_entries_2_valid_3 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_2_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3299) begin
          if (sectored_entries_2_data_3[0]) begin
            sectored_entries_2_valid_3 <= 1'h0;
          end else if (_T_739) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_2_valid_3 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1539) begin
                    sectored_entries_2_valid_3 <= _GEN_132;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1539) begin
                  sectored_entries_2_valid_3 <= _GEN_132;
                end
              end
            end
          end
        end else if (_T_739) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_2_valid_3 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1539) begin
                  sectored_entries_2_valid_3 <= _GEN_132;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1539) begin
                sectored_entries_2_valid_3 <= _GEN_132;
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_3 <= _GEN_715;
      end
    end else begin
      sectored_entries_2_valid_3 <= _GEN_496;
    end
    if (metaReset) begin
      sectored_entries_3_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1556) begin
            sectored_entries_3_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_3_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1556) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_0 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_3_data_1 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1556) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_1 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_3_data_2 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1556) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_2 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_3_data_3 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1556) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_3 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_3_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_3_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3470) begin
          if (sectored_entries_3_data_0[0]) begin
            sectored_entries_3_valid_0 <= 1'h0;
          end else if (_T_745) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_3_valid_0 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1556) begin
                    sectored_entries_3_valid_0 <= _GEN_151;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1556) begin
                  sectored_entries_3_valid_0 <= _GEN_151;
                end
              end
            end
          end
        end else if (_T_745) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_3_valid_0 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1556) begin
                  sectored_entries_3_valid_0 <= _GEN_151;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1556) begin
                sectored_entries_3_valid_0 <= _GEN_151;
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_0 <= _GEN_740;
      end
    end else begin
      sectored_entries_3_valid_0 <= _GEN_503;
    end
    if (metaReset) begin
      sectored_entries_3_valid_1 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_3_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3470) begin
          if (sectored_entries_3_data_1[0]) begin
            sectored_entries_3_valid_1 <= 1'h0;
          end else if (_T_745) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_3_valid_1 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1556) begin
                    sectored_entries_3_valid_1 <= _GEN_152;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1556) begin
                  sectored_entries_3_valid_1 <= _GEN_152;
                end
              end
            end
          end
        end else if (_T_745) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_3_valid_1 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1556) begin
                  sectored_entries_3_valid_1 <= _GEN_152;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1556) begin
                sectored_entries_3_valid_1 <= _GEN_152;
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_1 <= _GEN_741;
      end
    end else begin
      sectored_entries_3_valid_1 <= _GEN_504;
    end
    if (metaReset) begin
      sectored_entries_3_valid_2 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_3_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3470) begin
          if (sectored_entries_3_data_2[0]) begin
            sectored_entries_3_valid_2 <= 1'h0;
          end else if (_T_745) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_3_valid_2 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1556) begin
                    sectored_entries_3_valid_2 <= _GEN_153;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1556) begin
                  sectored_entries_3_valid_2 <= _GEN_153;
                end
              end
            end
          end
        end else if (_T_745) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_3_valid_2 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1556) begin
                  sectored_entries_3_valid_2 <= _GEN_153;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1556) begin
                sectored_entries_3_valid_2 <= _GEN_153;
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_2 <= _GEN_742;
      end
    end else begin
      sectored_entries_3_valid_2 <= _GEN_505;
    end
    if (metaReset) begin
      sectored_entries_3_valid_3 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_3_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3470) begin
          if (sectored_entries_3_data_3[0]) begin
            sectored_entries_3_valid_3 <= 1'h0;
          end else if (_T_745) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_3_valid_3 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1556) begin
                    sectored_entries_3_valid_3 <= _GEN_154;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1556) begin
                  sectored_entries_3_valid_3 <= _GEN_154;
                end
              end
            end
          end
        end else if (_T_745) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_3_valid_3 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1556) begin
                  sectored_entries_3_valid_3 <= _GEN_154;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1556) begin
                sectored_entries_3_valid_3 <= _GEN_154;
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_3 <= _GEN_743;
      end
    end else begin
      sectored_entries_3_valid_3 <= _GEN_506;
    end
    if (metaReset) begin
      sectored_entries_4_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1573) begin
            sectored_entries_4_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_4_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1573) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_0 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_4_data_1 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1573) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_1 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_4_data_2 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1573) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_2 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_4_data_3 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1573) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_3 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_4_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_4_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3641) begin
          if (sectored_entries_4_data_0[0]) begin
            sectored_entries_4_valid_0 <= 1'h0;
          end else if (_T_751) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_4_valid_0 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1573) begin
                    sectored_entries_4_valid_0 <= _GEN_173;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1573) begin
                  sectored_entries_4_valid_0 <= _GEN_173;
                end
              end
            end
          end
        end else if (_T_751) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_4_valid_0 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1573) begin
                  sectored_entries_4_valid_0 <= _GEN_173;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1573) begin
                sectored_entries_4_valid_0 <= _GEN_173;
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_0 <= _GEN_768;
      end
    end else begin
      sectored_entries_4_valid_0 <= _GEN_513;
    end
    if (metaReset) begin
      sectored_entries_4_valid_1 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_4_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3641) begin
          if (sectored_entries_4_data_1[0]) begin
            sectored_entries_4_valid_1 <= 1'h0;
          end else if (_T_751) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_4_valid_1 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1573) begin
                    sectored_entries_4_valid_1 <= _GEN_174;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1573) begin
                  sectored_entries_4_valid_1 <= _GEN_174;
                end
              end
            end
          end
        end else if (_T_751) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_4_valid_1 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1573) begin
                  sectored_entries_4_valid_1 <= _GEN_174;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1573) begin
                sectored_entries_4_valid_1 <= _GEN_174;
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_1 <= _GEN_769;
      end
    end else begin
      sectored_entries_4_valid_1 <= _GEN_514;
    end
    if (metaReset) begin
      sectored_entries_4_valid_2 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_4_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3641) begin
          if (sectored_entries_4_data_2[0]) begin
            sectored_entries_4_valid_2 <= 1'h0;
          end else if (_T_751) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_4_valid_2 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1573) begin
                    sectored_entries_4_valid_2 <= _GEN_175;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1573) begin
                  sectored_entries_4_valid_2 <= _GEN_175;
                end
              end
            end
          end
        end else if (_T_751) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_4_valid_2 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1573) begin
                  sectored_entries_4_valid_2 <= _GEN_175;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1573) begin
                sectored_entries_4_valid_2 <= _GEN_175;
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_2 <= _GEN_770;
      end
    end else begin
      sectored_entries_4_valid_2 <= _GEN_515;
    end
    if (metaReset) begin
      sectored_entries_4_valid_3 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_4_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3641) begin
          if (sectored_entries_4_data_3[0]) begin
            sectored_entries_4_valid_3 <= 1'h0;
          end else if (_T_751) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_4_valid_3 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1573) begin
                    sectored_entries_4_valid_3 <= _GEN_176;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1573) begin
                  sectored_entries_4_valid_3 <= _GEN_176;
                end
              end
            end
          end
        end else if (_T_751) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_4_valid_3 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1573) begin
                  sectored_entries_4_valid_3 <= _GEN_176;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1573) begin
                sectored_entries_4_valid_3 <= _GEN_176;
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_3 <= _GEN_771;
      end
    end else begin
      sectored_entries_4_valid_3 <= _GEN_516;
    end
    if (metaReset) begin
      sectored_entries_5_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1590) begin
            sectored_entries_5_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_5_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1590) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_0 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_5_data_1 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1590) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_1 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_5_data_2 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1590) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_2 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_5_data_3 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1590) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_3 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_5_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_5_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3812) begin
          if (sectored_entries_5_data_0[0]) begin
            sectored_entries_5_valid_0 <= 1'h0;
          end else if (_T_757) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_5_valid_0 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1590) begin
                    sectored_entries_5_valid_0 <= _GEN_195;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1590) begin
                  sectored_entries_5_valid_0 <= _GEN_195;
                end
              end
            end
          end
        end else if (_T_757) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_5_valid_0 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1590) begin
                  sectored_entries_5_valid_0 <= _GEN_195;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1590) begin
                sectored_entries_5_valid_0 <= _GEN_195;
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_0 <= _GEN_796;
      end
    end else begin
      sectored_entries_5_valid_0 <= _GEN_523;
    end
    if (metaReset) begin
      sectored_entries_5_valid_1 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_5_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3812) begin
          if (sectored_entries_5_data_1[0]) begin
            sectored_entries_5_valid_1 <= 1'h0;
          end else if (_T_757) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_5_valid_1 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1590) begin
                    sectored_entries_5_valid_1 <= _GEN_196;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1590) begin
                  sectored_entries_5_valid_1 <= _GEN_196;
                end
              end
            end
          end
        end else if (_T_757) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_5_valid_1 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1590) begin
                  sectored_entries_5_valid_1 <= _GEN_196;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1590) begin
                sectored_entries_5_valid_1 <= _GEN_196;
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_1 <= _GEN_797;
      end
    end else begin
      sectored_entries_5_valid_1 <= _GEN_524;
    end
    if (metaReset) begin
      sectored_entries_5_valid_2 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_5_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3812) begin
          if (sectored_entries_5_data_2[0]) begin
            sectored_entries_5_valid_2 <= 1'h0;
          end else if (_T_757) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_5_valid_2 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1590) begin
                    sectored_entries_5_valid_2 <= _GEN_197;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1590) begin
                  sectored_entries_5_valid_2 <= _GEN_197;
                end
              end
            end
          end
        end else if (_T_757) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_5_valid_2 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1590) begin
                  sectored_entries_5_valid_2 <= _GEN_197;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1590) begin
                sectored_entries_5_valid_2 <= _GEN_197;
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_2 <= _GEN_798;
      end
    end else begin
      sectored_entries_5_valid_2 <= _GEN_525;
    end
    if (metaReset) begin
      sectored_entries_5_valid_3 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_5_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3812) begin
          if (sectored_entries_5_data_3[0]) begin
            sectored_entries_5_valid_3 <= 1'h0;
          end else if (_T_757) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_5_valid_3 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1590) begin
                    sectored_entries_5_valid_3 <= _GEN_198;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1590) begin
                  sectored_entries_5_valid_3 <= _GEN_198;
                end
              end
            end
          end
        end else if (_T_757) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_5_valid_3 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1590) begin
                  sectored_entries_5_valid_3 <= _GEN_198;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1590) begin
                sectored_entries_5_valid_3 <= _GEN_198;
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_3 <= _GEN_799;
      end
    end else begin
      sectored_entries_5_valid_3 <= _GEN_526;
    end
    if (metaReset) begin
      sectored_entries_6_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1607) begin
            sectored_entries_6_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_6_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1607) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_0 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_6_data_1 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1607) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_1 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_6_data_2 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1607) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_2 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_6_data_3 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1607) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_3 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_6_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_6_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3983) begin
          if (sectored_entries_6_data_0[0]) begin
            sectored_entries_6_valid_0 <= 1'h0;
          end else if (_T_763) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_6_valid_0 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1607) begin
                    sectored_entries_6_valid_0 <= _GEN_217;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1607) begin
                  sectored_entries_6_valid_0 <= _GEN_217;
                end
              end
            end
          end
        end else if (_T_763) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_6_valid_0 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1607) begin
                  sectored_entries_6_valid_0 <= _GEN_217;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1607) begin
                sectored_entries_6_valid_0 <= _GEN_217;
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_0 <= _GEN_824;
      end
    end else begin
      sectored_entries_6_valid_0 <= _GEN_533;
    end
    if (metaReset) begin
      sectored_entries_6_valid_1 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_6_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3983) begin
          if (sectored_entries_6_data_1[0]) begin
            sectored_entries_6_valid_1 <= 1'h0;
          end else if (_T_763) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_6_valid_1 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1607) begin
                    sectored_entries_6_valid_1 <= _GEN_218;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1607) begin
                  sectored_entries_6_valid_1 <= _GEN_218;
                end
              end
            end
          end
        end else if (_T_763) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_6_valid_1 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1607) begin
                  sectored_entries_6_valid_1 <= _GEN_218;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1607) begin
                sectored_entries_6_valid_1 <= _GEN_218;
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_1 <= _GEN_825;
      end
    end else begin
      sectored_entries_6_valid_1 <= _GEN_534;
    end
    if (metaReset) begin
      sectored_entries_6_valid_2 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_6_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3983) begin
          if (sectored_entries_6_data_2[0]) begin
            sectored_entries_6_valid_2 <= 1'h0;
          end else if (_T_763) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_6_valid_2 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1607) begin
                    sectored_entries_6_valid_2 <= _GEN_219;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1607) begin
                  sectored_entries_6_valid_2 <= _GEN_219;
                end
              end
            end
          end
        end else if (_T_763) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_6_valid_2 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1607) begin
                  sectored_entries_6_valid_2 <= _GEN_219;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1607) begin
                sectored_entries_6_valid_2 <= _GEN_219;
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_2 <= _GEN_826;
      end
    end else begin
      sectored_entries_6_valid_2 <= _GEN_535;
    end
    if (metaReset) begin
      sectored_entries_6_valid_3 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_6_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3983) begin
          if (sectored_entries_6_data_3[0]) begin
            sectored_entries_6_valid_3 <= 1'h0;
          end else if (_T_763) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_6_valid_3 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1607) begin
                    sectored_entries_6_valid_3 <= _GEN_220;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1607) begin
                  sectored_entries_6_valid_3 <= _GEN_220;
                end
              end
            end
          end
        end else if (_T_763) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_6_valid_3 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1607) begin
                  sectored_entries_6_valid_3 <= _GEN_220;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1607) begin
                sectored_entries_6_valid_3 <= _GEN_220;
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_3 <= _GEN_827;
      end
    end else begin
      sectored_entries_6_valid_3 <= _GEN_536;
    end
    if (metaReset) begin
      sectored_entries_7_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1624) begin
            sectored_entries_7_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_7_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1624) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_0 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_7_data_1 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1624) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_1 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_7_data_2 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1624) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_2 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_7_data_3 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1624) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_3 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_7_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_7_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_4154) begin
          if (sectored_entries_7_data_0[0]) begin
            sectored_entries_7_valid_0 <= 1'h0;
          end else if (_T_769) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_7_valid_0 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1624) begin
                    sectored_entries_7_valid_0 <= _GEN_239;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1624) begin
                  sectored_entries_7_valid_0 <= _GEN_239;
                end
              end
            end
          end
        end else if (_T_769) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_7_valid_0 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1624) begin
                  sectored_entries_7_valid_0 <= _GEN_239;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1624) begin
                sectored_entries_7_valid_0 <= _GEN_239;
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_0 <= _GEN_852;
      end
    end else begin
      sectored_entries_7_valid_0 <= _GEN_543;
    end
    if (metaReset) begin
      sectored_entries_7_valid_1 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_7_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_4154) begin
          if (sectored_entries_7_data_1[0]) begin
            sectored_entries_7_valid_1 <= 1'h0;
          end else if (_T_769) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_7_valid_1 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1624) begin
                    sectored_entries_7_valid_1 <= _GEN_240;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1624) begin
                  sectored_entries_7_valid_1 <= _GEN_240;
                end
              end
            end
          end
        end else if (_T_769) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_7_valid_1 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1624) begin
                  sectored_entries_7_valid_1 <= _GEN_240;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1624) begin
                sectored_entries_7_valid_1 <= _GEN_240;
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_1 <= _GEN_853;
      end
    end else begin
      sectored_entries_7_valid_1 <= _GEN_544;
    end
    if (metaReset) begin
      sectored_entries_7_valid_2 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_7_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_4154) begin
          if (sectored_entries_7_data_2[0]) begin
            sectored_entries_7_valid_2 <= 1'h0;
          end else if (_T_769) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_7_valid_2 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1624) begin
                    sectored_entries_7_valid_2 <= _GEN_241;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1624) begin
                  sectored_entries_7_valid_2 <= _GEN_241;
                end
              end
            end
          end
        end else if (_T_769) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_7_valid_2 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1624) begin
                  sectored_entries_7_valid_2 <= _GEN_241;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1624) begin
                sectored_entries_7_valid_2 <= _GEN_241;
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_2 <= _GEN_854;
      end
    end else begin
      sectored_entries_7_valid_2 <= _GEN_545;
    end
    if (metaReset) begin
      sectored_entries_7_valid_3 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_7_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_4154) begin
          if (sectored_entries_7_data_3[0]) begin
            sectored_entries_7_valid_3 <= 1'h0;
          end else if (_T_769) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_7_valid_3 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1624) begin
                    sectored_entries_7_valid_3 <= _GEN_242;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1624) begin
                  sectored_entries_7_valid_3 <= _GEN_242;
                end
              end
            end
          end
        end else if (_T_769) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_7_valid_3 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1624) begin
                  sectored_entries_7_valid_3 <= _GEN_242;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1624) begin
                sectored_entries_7_valid_3 <= _GEN_242;
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_3 <= _GEN_855;
      end
    end else begin
      sectored_entries_7_valid_3 <= _GEN_546;
    end
    if (metaReset) begin
      superpage_entries_0_level <= 2'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1440) begin
            superpage_entries_0_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_0_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1440) begin
            superpage_entries_0_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_0_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1440) begin
            superpage_entries_0_data_0 <= _T_1438;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_0_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      superpage_entries_0_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_0) begin
          superpage_entries_0_valid_0 <= 1'h0;
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_1439) begin
              superpage_entries_0_valid_0 <= _GEN_67;
            end
          end
        end
      end else begin
        superpage_entries_0_valid_0 <= _GEN_862;
      end
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          superpage_entries_0_valid_0 <= _GEN_67;
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_level <= 2'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1456) begin
            superpage_entries_1_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1456) begin
            superpage_entries_1_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1456) begin
            superpage_entries_1_data_0 <= _T_1438;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      superpage_entries_1_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_1) begin
          superpage_entries_1_valid_0 <= 1'h0;
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_1439) begin
              superpage_entries_1_valid_0 <= _GEN_71;
            end
          end
        end
      end else begin
        superpage_entries_1_valid_0 <= _GEN_866;
      end
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          superpage_entries_1_valid_0 <= _GEN_71;
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_level <= 2'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1472) begin
            superpage_entries_2_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1472) begin
            superpage_entries_2_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1472) begin
            superpage_entries_2_data_0 <= _T_1438;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      superpage_entries_2_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_2) begin
          superpage_entries_2_valid_0 <= 1'h0;
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_1439) begin
              superpage_entries_2_valid_0 <= _GEN_75;
            end
          end
        end
      end else begin
        superpage_entries_2_valid_0 <= _GEN_870;
      end
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          superpage_entries_2_valid_0 <= _GEN_75;
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_level <= 2'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1488) begin
            superpage_entries_3_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1488) begin
            superpage_entries_3_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1488) begin
            superpage_entries_3_data_0 <= _T_1438;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      superpage_entries_3_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_3) begin
          superpage_entries_3_valid_0 <= 1'h0;
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_1439) begin
              superpage_entries_3_valid_0 <= _GEN_79;
            end
          end
        end
      end else begin
        superpage_entries_3_valid_0 <= _GEN_874;
      end
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          superpage_entries_3_valid_0 <= _GEN_79;
        end
      end
    end
    if (metaReset) begin
      special_entry_level <= 2'h0;
    end else if (_T_1385) begin
      if (~io_ptw_resp_bits_homogeneous) begin
        special_entry_level <= io_ptw_resp_bits_level;
      end
    end
    if (metaReset) begin
      special_entry_tag <= 27'h0;
    end else if (_T_1385) begin
      if (~io_ptw_resp_bits_homogeneous) begin
        special_entry_tag <= r_refill_tag;
      end
    end
    if (metaReset) begin
      special_entry_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (~io_ptw_resp_bits_homogeneous) begin
        special_entry_data_0 <= _T_1438;
      end
    end
    if (metaReset) begin
      special_entry_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      special_entry_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_994) begin
          special_entry_valid_0 <= 1'h0;
        end else if (_T_1385) begin
          special_entry_valid_0 <= _GEN_355;
        end
      end else begin
        special_entry_valid_0 <= _GEN_878;
      end
    end else if (_T_1385) begin
      special_entry_valid_0 <= _GEN_355;
    end
    if (metaReset) begin
      state <= 2'h0;
    end else if (reset) begin
      state <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      state <= 2'h0;
    end else if (_T_2941) begin
      state <= 2'h3;
    end else if (io_ptw_resp_valid) begin
      state <= 2'h0;
    end else if (_T_2941) begin
      state <= 2'h3;
    end else if (_T_324) begin
      if (io_ptw_req_ready) begin
        if (io_sfence_valid) begin
          state <= 2'h3;
        end else begin
          state <= 2'h2;
        end
      end else if (io_sfence_valid) begin
        state <= 2'h0;
      end else if (_T_2809) begin
        state <= 2'h1;
      end
    end else if (_T_2809) begin
      state <= 2'h1;
    end
    if (metaReset) begin
      r_refill_tag <= 27'h0;
    end else if (_T_2809) begin
      r_refill_tag <= vpn;
    end
    if (metaReset) begin
      r_superpage_repl_addr <= 2'h0;
    end else if (_T_2809) begin
      if (_T_2830) begin
        r_superpage_repl_addr <= _T_2824[1:0];
      end else if (_T_2832) begin
        r_superpage_repl_addr <= 2'h0;
      end else if (_T_2833) begin
        r_superpage_repl_addr <= 2'h1;
      end else if (_T_2834) begin
        r_superpage_repl_addr <= 2'h2;
      end else begin
        r_superpage_repl_addr <= 2'h3;
      end
    end
    if (metaReset) begin
      r_sectored_repl_addr <= 3'h0;
    end else if (_T_2809) begin
      if (_T_2895) begin
        r_sectored_repl_addr <= _T_2861[2:0];
      end else if (_T_2897) begin
        r_sectored_repl_addr <= 3'h0;
      end else if (_T_2898) begin
        r_sectored_repl_addr <= 3'h1;
      end else if (_T_2899) begin
        r_sectored_repl_addr <= 3'h2;
      end else if (_T_2900) begin
        r_sectored_repl_addr <= 3'h3;
      end else if (_T_2901) begin
        r_sectored_repl_addr <= 3'h4;
      end else if (_T_2902) begin
        r_sectored_repl_addr <= 3'h5;
      end else if (_T_2903) begin
        r_sectored_repl_addr <= 3'h6;
      end else begin
        r_sectored_repl_addr <= 3'h7;
      end
    end
    if (metaReset) begin
      r_sectored_hit_addr <= 3'h0;
    end else if (_T_2809) begin
      r_sectored_hit_addr <= _T_2582;
    end
    if (metaReset) begin
      r_sectored_hit <= 1'h0;
    end else if (_T_2809) begin
      r_sectored_hit <= _T_2564;
    end
    if (metaReset) begin
      vpoffset_cfg_value <= 27'h0;
    end else if (reset) begin
      vpoffset_cfg_value <= 27'h0;
    end else begin
      vpoffset_cfg_value <= io_ptw_vpoffset_bits_value;
    end
    if (metaReset) begin
      requestedVPN <= 27'h0;
    end else if (io_ptw_req_bits_valid) begin
      requestedVPN <= io_ptw_req_bits_bits_addr;
    end
    if (metaReset) begin
      _T_2554 <= 7'h0;
    end else if (_T_2557) begin
      if (_T_2564) begin
        _T_2554 <= _T_2609[7:1];
      end
    end
    if (metaReset) begin
      _T_2556 <= 3'h0;
    end else if (_T_2557) begin
      if (_T_2614) begin
        _T_2556 <= _T_2641[3:1];
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_sfence_valid & ~_T_2949) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TLB.scala:414 assert(!io.sfence.bits.rs1 || (io.sfence.bits.addr >> pgIdxBits) === vpn)\n"); // @[TLB.scala 414:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_sfence_valid & ~_T_2949) begin
          $fatal; // @[TLB.scala 414:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    TLB_state <= TLB_xor0;
    if (!(TLB_cov_read_data)) begin
      TLB_covSum <= TLB_covSum + 1'h1;
    end
    if (metaReset) begin
      TLB_metaAssert <= 1'h0;
    end else begin
      TLB_metaAssert <= TLB_metaAssert | TLB_or0;
    end
  end
  always @(posedge clock) begin
    if(TLB_cov_write_en & TLB_cov_write_mask) begin
      TLB_cov[TLB_cov_write_addr] <= TLB_cov_write_data; // @[Coverage map for TLB]
    end
  end
endmodule
module AMOALU(
  input  [7:0]  io_mask,
  input  [4:0]  io_cmd,
  input  [63:0] io_lhs,
  input  [63:0] io_rhs,
  output [63:0] io_out,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  _T_10; // @[AMOALU.scala 64:20]
  wire  _T_11; // @[AMOALU.scala 64:43]
  wire  max; // @[AMOALU.scala 64:33]
  wire  _T_12; // @[AMOALU.scala 65:20]
  wire  _T_13; // @[AMOALU.scala 65:43]
  wire  min; // @[AMOALU.scala 65:33]
  wire  add; // @[AMOALU.scala 66:20]
  wire  _T_14; // @[AMOALU.scala 67:26]
  wire  _T_15; // @[AMOALU.scala 67:48]
  wire  logic_and; // @[AMOALU.scala 67:38]
  wire  _T_16; // @[AMOALU.scala 68:26]
  wire  logic_xor; // @[AMOALU.scala 68:39]
  wire [31:0] _T_20; // @[AMOALU.scala 72:79]
  wire [63:0] _T_21; // @[AMOALU.scala 72:98]
  wire [63:0] _T_23; // @[AMOALU.scala 73:13]
  wire [63:0] _T_24; // @[AMOALU.scala 73:31]
  wire [63:0] adder_out; // @[AMOALU.scala 73:21]
  wire [4:0] _T_28; // @[AMOALU.scala 86:17]
  wire  _T_30; // @[AMOALU.scala 86:25]
  wire  _T_33; // @[AMOALU.scala 88:18]
  wire  _T_36; // @[AMOALU.scala 80:24]
  wire  _T_39; // @[AMOALU.scala 80:53]
  wire  _T_42; // @[AMOALU.scala 79:35]
  wire  _T_43; // @[AMOALU.scala 80:69]
  wire  _T_44; // @[AMOALU.scala 80:38]
  wire  _T_47; // @[AMOALU.scala 88:58]
  wire  _T_48; // @[AMOALU.scala 88:10]
  wire  _T_56; // @[AMOALU.scala 88:18]
  wire  _T_62; // @[AMOALU.scala 88:58]
  wire  _T_63; // @[AMOALU.scala 88:10]
  wire  less; // @[Mux.scala 31:69]
  wire  _T_64; // @[AMOALU.scala 94:23]
  wire [63:0] minmax; // @[AMOALU.scala 94:19]
  wire [63:0] _T_65; // @[AMOALU.scala 96:27]
  wire [63:0] _T_66; // @[AMOALU.scala 96:8]
  wire [63:0] _T_67; // @[AMOALU.scala 97:27]
  wire [63:0] _T_68; // @[AMOALU.scala 97:8]
  wire [63:0] logic_; // @[AMOALU.scala 96:42]
  wire  _T_69; // @[AMOALU.scala 100:19]
  wire [63:0] _T_70; // @[AMOALU.scala 100:8]
  wire [63:0] out; // @[AMOALU.scala 99:8]
  wire [7:0] _T_80; // @[Bitwise.scala 72:12]
  wire [7:0] _T_82; // @[Bitwise.scala 72:12]
  wire [7:0] _T_84; // @[Bitwise.scala 72:12]
  wire [7:0] _T_86; // @[Bitwise.scala 72:12]
  wire [7:0] _T_88; // @[Bitwise.scala 72:12]
  wire [7:0] _T_90; // @[Bitwise.scala 72:12]
  wire [7:0] _T_92; // @[Bitwise.scala 72:12]
  wire [7:0] _T_94; // @[Bitwise.scala 72:12]
  wire [63:0] wmask; // @[Cat.scala 30:58]
  wire [63:0] _T_101; // @[AMOALU.scala 104:19]
  wire [63:0] _T_103; // @[AMOALU.scala 104:34]
  wire [29:0] AMOALU_covSum;
  assign _T_10 = io_cmd == 5'hd; // @[AMOALU.scala 64:20]
  assign _T_11 = io_cmd == 5'hf; // @[AMOALU.scala 64:43]
  assign max = _T_10 | _T_11; // @[AMOALU.scala 64:33]
  assign _T_12 = io_cmd == 5'hc; // @[AMOALU.scala 65:20]
  assign _T_13 = io_cmd == 5'he; // @[AMOALU.scala 65:43]
  assign min = _T_12 | _T_13; // @[AMOALU.scala 65:33]
  assign add = io_cmd == 5'h8; // @[AMOALU.scala 66:20]
  assign _T_14 = io_cmd == 5'ha; // @[AMOALU.scala 67:26]
  assign _T_15 = io_cmd == 5'hb; // @[AMOALU.scala 67:48]
  assign logic_and = _T_14 | _T_15; // @[AMOALU.scala 67:38]
  assign _T_16 = io_cmd == 5'h9; // @[AMOALU.scala 68:26]
  assign logic_xor = _T_16 | _T_14; // @[AMOALU.scala 68:39]
  assign _T_20 = {~io_mask[3], 31'h0}; // @[AMOALU.scala 72:79]
  assign _T_21 = {{32'd0}, _T_20}; // @[AMOALU.scala 72:98]
  assign _T_23 = io_lhs & ~_T_21; // @[AMOALU.scala 73:13]
  assign _T_24 = io_rhs & ~_T_21; // @[AMOALU.scala 73:31]
  assign adder_out = _T_23 + _T_24; // @[AMOALU.scala 73:21]
  assign _T_28 = io_cmd & 5'h2; // @[AMOALU.scala 86:17]
  assign _T_30 = _T_28 == 5'h0; // @[AMOALU.scala 86:25]
  assign _T_33 = io_lhs[63] == io_rhs[63]; // @[AMOALU.scala 88:18]
  assign _T_36 = io_lhs[63:32] < io_rhs[63:32]; // @[AMOALU.scala 80:24]
  assign _T_39 = io_lhs[63:32] == io_rhs[63:32]; // @[AMOALU.scala 80:53]
  assign _T_42 = io_lhs[31:0] < io_rhs[31:0]; // @[AMOALU.scala 79:35]
  assign _T_43 = _T_39 & _T_42; // @[AMOALU.scala 80:69]
  assign _T_44 = _T_36 | _T_43; // @[AMOALU.scala 80:38]
  assign _T_47 = _T_30 ? io_lhs[63] : io_rhs[63]; // @[AMOALU.scala 88:58]
  assign _T_48 = _T_33 ? _T_44 : _T_47; // @[AMOALU.scala 88:10]
  assign _T_56 = io_lhs[31] == io_rhs[31]; // @[AMOALU.scala 88:18]
  assign _T_62 = _T_30 ? io_lhs[31] : io_rhs[31]; // @[AMOALU.scala 88:58]
  assign _T_63 = _T_56 ? _T_42 : _T_62; // @[AMOALU.scala 88:10]
  assign less = io_mask[4] ? _T_48 : _T_63; // @[Mux.scala 31:69]
  assign _T_64 = less ? min : max; // @[AMOALU.scala 94:23]
  assign minmax = _T_64 ? io_lhs : io_rhs; // @[AMOALU.scala 94:19]
  assign _T_65 = io_lhs & io_rhs; // @[AMOALU.scala 96:27]
  assign _T_66 = logic_and ? _T_65 : 64'h0; // @[AMOALU.scala 96:8]
  assign _T_67 = io_lhs ^ io_rhs; // @[AMOALU.scala 97:27]
  assign _T_68 = logic_xor ? _T_67 : 64'h0; // @[AMOALU.scala 97:8]
  assign logic_ = _T_66 | _T_68; // @[AMOALU.scala 96:42]
  assign _T_69 = logic_and | logic_xor; // @[AMOALU.scala 100:19]
  assign _T_70 = _T_69 ? logic_ : minmax; // @[AMOALU.scala 100:8]
  assign out = add ? adder_out : _T_70; // @[AMOALU.scala 99:8]
  assign _T_80 = io_mask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_82 = io_mask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_84 = io_mask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_86 = io_mask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_88 = io_mask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_90 = io_mask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_92 = io_mask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_94 = io_mask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign wmask = {_T_94,_T_92,_T_90,_T_88,_T_86,_T_84,_T_82,_T_80}; // @[Cat.scala 30:58]
  assign _T_101 = wmask & out; // @[AMOALU.scala 104:19]
  assign _T_103 = ~wmask & io_lhs; // @[AMOALU.scala 104:34]
  assign io_out = _T_101 | _T_103; // @[AMOALU.scala 104:10]
  assign AMOALU_covSum = 30'h0;
  assign io_covSum = AMOALU_covSum;
  assign metaAssert = 1'h0;
endmodule
module ICache(
  input         clock,
  input         reset,
  input         auto_master_out_a_ready,
  output        auto_master_out_a_valid,
  output [31:0] auto_master_out_a_bits_address,
  input         auto_master_out_d_valid,
  input  [2:0]  auto_master_out_d_bits_opcode,
  input  [3:0]  auto_master_out_d_bits_size,
  input  [63:0] auto_master_out_d_bits_data,
  input         auto_master_out_d_bits_corrupt,
  output        io_req_ready,
  input         io_req_valid,
  input  [38:0] io_req_bits_addr,
  input  [31:0] io_s1_paddr,
  input         io_s1_kill,
  input         io_s2_kill,
  output        io_resp_valid,
  output [31:0] io_resp_bits_data,
  output        io_resp_bits_ae,
  input         io_invalidate,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [20:0] tag_array_0 [0:63]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_0;
  wire [20:0] tag_array_0_tag_rdata_data; // @[DescribedSRAM.scala 23:21]
  wire [5:0] tag_array_0_tag_rdata_addr; // @[DescribedSRAM.scala 23:21]
  wire [20:0] tag_array_0__T_256_data; // @[DescribedSRAM.scala 23:21]
  wire [5:0] tag_array_0__T_256_addr; // @[DescribedSRAM.scala 23:21]
  wire  tag_array_0__T_256_mask; // @[DescribedSRAM.scala 23:21]
  wire  tag_array_0__T_256_en; // @[DescribedSRAM.scala 23:21]
  reg  tag_array_0_tag_rdata_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [5:0] tag_array_0_tag_rdata_addr_pipe_0;
  reg [31:0] _RAND_2;
  reg [20:0] tag_array_1 [0:63]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_3;
  wire [20:0] tag_array_1_tag_rdata_data; // @[DescribedSRAM.scala 23:21]
  wire [5:0] tag_array_1_tag_rdata_addr; // @[DescribedSRAM.scala 23:21]
  wire [20:0] tag_array_1__T_256_data; // @[DescribedSRAM.scala 23:21]
  wire [5:0] tag_array_1__T_256_addr; // @[DescribedSRAM.scala 23:21]
  wire  tag_array_1__T_256_mask; // @[DescribedSRAM.scala 23:21]
  wire  tag_array_1__T_256_en; // @[DescribedSRAM.scala 23:21]
  reg  tag_array_1_tag_rdata_en_pipe_0;
  reg [31:0] _RAND_4;
  reg [5:0] tag_array_1_tag_rdata_addr_pipe_0;
  reg [31:0] _RAND_5;
  reg [20:0] tag_array_2 [0:63]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_6;
  wire [20:0] tag_array_2_tag_rdata_data; // @[DescribedSRAM.scala 23:21]
  wire [5:0] tag_array_2_tag_rdata_addr; // @[DescribedSRAM.scala 23:21]
  wire [20:0] tag_array_2__T_256_data; // @[DescribedSRAM.scala 23:21]
  wire [5:0] tag_array_2__T_256_addr; // @[DescribedSRAM.scala 23:21]
  wire  tag_array_2__T_256_mask; // @[DescribedSRAM.scala 23:21]
  wire  tag_array_2__T_256_en; // @[DescribedSRAM.scala 23:21]
  reg  tag_array_2_tag_rdata_en_pipe_0;
  reg [31:0] _RAND_7;
  reg [5:0] tag_array_2_tag_rdata_addr_pipe_0;
  reg [31:0] _RAND_8;
  reg [20:0] tag_array_3 [0:63]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_9;
  wire [20:0] tag_array_3_tag_rdata_data; // @[DescribedSRAM.scala 23:21]
  wire [5:0] tag_array_3_tag_rdata_addr; // @[DescribedSRAM.scala 23:21]
  wire [20:0] tag_array_3__T_256_data; // @[DescribedSRAM.scala 23:21]
  wire [5:0] tag_array_3__T_256_addr; // @[DescribedSRAM.scala 23:21]
  wire  tag_array_3__T_256_mask; // @[DescribedSRAM.scala 23:21]
  wire  tag_array_3__T_256_en; // @[DescribedSRAM.scala 23:21]
  reg  tag_array_3_tag_rdata_en_pipe_0;
  reg [31:0] _RAND_10;
  reg [5:0] tag_array_3_tag_rdata_addr_pipe_0;
  reg [31:0] _RAND_11;
  reg [31:0] data_arrays_0_0 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_12;
  wire [31:0] data_arrays_0_0__T_513_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_0__T_513_addr; // @[DescribedSRAM.scala 23:21]
  wire [31:0] data_arrays_0_0__T_495_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_0__T_495_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_0__T_495_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_0__T_495_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_0__T_513_en_pipe_0;
  reg [31:0] _RAND_13;
  reg [8:0] data_arrays_0_0__T_513_addr_pipe_0;
  reg [31:0] _RAND_14;
  reg [31:0] data_arrays_0_1 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_15;
  wire [31:0] data_arrays_0_1__T_513_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_1__T_513_addr; // @[DescribedSRAM.scala 23:21]
  wire [31:0] data_arrays_0_1__T_495_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_1__T_495_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_1__T_495_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_1__T_495_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_1__T_513_en_pipe_0;
  reg [31:0] _RAND_16;
  reg [8:0] data_arrays_0_1__T_513_addr_pipe_0;
  reg [31:0] _RAND_17;
  reg [31:0] data_arrays_0_2 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_18;
  wire [31:0] data_arrays_0_2__T_513_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_2__T_513_addr; // @[DescribedSRAM.scala 23:21]
  wire [31:0] data_arrays_0_2__T_495_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_2__T_495_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_2__T_495_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_2__T_495_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_2__T_513_en_pipe_0;
  reg [31:0] _RAND_19;
  reg [8:0] data_arrays_0_2__T_513_addr_pipe_0;
  reg [31:0] _RAND_20;
  reg [31:0] data_arrays_0_3 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_21;
  wire [31:0] data_arrays_0_3__T_513_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_3__T_513_addr; // @[DescribedSRAM.scala 23:21]
  wire [31:0] data_arrays_0_3__T_495_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_0_3__T_495_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_3__T_495_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_0_3__T_495_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_0_3__T_513_en_pipe_0;
  reg [31:0] _RAND_22;
  reg [8:0] data_arrays_0_3__T_513_addr_pipe_0;
  reg [31:0] _RAND_23;
  reg [31:0] data_arrays_1_0 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_24;
  wire [31:0] data_arrays_1_0__T_583_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_1_0__T_583_addr; // @[DescribedSRAM.scala 23:21]
  wire [31:0] data_arrays_1_0__T_565_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_1_0__T_565_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_1_0__T_565_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_1_0__T_565_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_1_0__T_583_en_pipe_0;
  reg [31:0] _RAND_25;
  reg [8:0] data_arrays_1_0__T_583_addr_pipe_0;
  reg [31:0] _RAND_26;
  reg [31:0] data_arrays_1_1 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_27;
  wire [31:0] data_arrays_1_1__T_583_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_1_1__T_583_addr; // @[DescribedSRAM.scala 23:21]
  wire [31:0] data_arrays_1_1__T_565_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_1_1__T_565_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_1_1__T_565_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_1_1__T_565_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_1_1__T_583_en_pipe_0;
  reg [31:0] _RAND_28;
  reg [8:0] data_arrays_1_1__T_583_addr_pipe_0;
  reg [31:0] _RAND_29;
  reg [31:0] data_arrays_1_2 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_30;
  wire [31:0] data_arrays_1_2__T_583_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_1_2__T_583_addr; // @[DescribedSRAM.scala 23:21]
  wire [31:0] data_arrays_1_2__T_565_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_1_2__T_565_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_1_2__T_565_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_1_2__T_565_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_1_2__T_583_en_pipe_0;
  reg [31:0] _RAND_31;
  reg [8:0] data_arrays_1_2__T_583_addr_pipe_0;
  reg [31:0] _RAND_32;
  reg [31:0] data_arrays_1_3 [0:511]; // @[DescribedSRAM.scala 23:21]
  reg [31:0] _RAND_33;
  wire [31:0] data_arrays_1_3__T_583_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_1_3__T_583_addr; // @[DescribedSRAM.scala 23:21]
  wire [31:0] data_arrays_1_3__T_565_data; // @[DescribedSRAM.scala 23:21]
  wire [8:0] data_arrays_1_3__T_565_addr; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_1_3__T_565_mask; // @[DescribedSRAM.scala 23:21]
  wire  data_arrays_1_3__T_565_en; // @[DescribedSRAM.scala 23:21]
  reg  data_arrays_1_3__T_583_en_pipe_0;
  reg [31:0] _RAND_34;
  reg [8:0] data_arrays_1_3__T_583_addr_pipe_0;
  reg [31:0] _RAND_35;
  reg  s1_valid; // @[ICache.scala 136:21]
  reg [31:0] _RAND_36;
  reg [255:0] vb_array; // @[ICache.scala 195:21]
  reg [255:0] _RAND_37;
  wire [6:0] _T_322; // @[Cat.scala 30:58]
  wire [255:0] _T_323; // @[ICache.scala 222:25]
  wire  _T_329; // @[ICache.scala 225:33]
  wire  s1_tag_hit_0; // @[ICache.scala 225:26]
  wire [6:0] _T_350; // @[Cat.scala 30:58]
  wire [255:0] _T_351; // @[ICache.scala 222:25]
  wire  _T_357; // @[ICache.scala 225:33]
  wire  s1_tag_hit_1; // @[ICache.scala 225:26]
  wire  _T_141; // @[ICache.scala 138:35]
  wire [7:0] _T_378; // @[Cat.scala 30:58]
  wire [255:0] _T_379; // @[ICache.scala 222:25]
  wire  _T_385; // @[ICache.scala 225:33]
  wire  s1_tag_hit_2; // @[ICache.scala 225:26]
  wire  _T_142; // @[ICache.scala 138:35]
  wire [7:0] _T_406; // @[Cat.scala 30:58]
  wire [255:0] _T_407; // @[ICache.scala 222:25]
  wire  _T_413; // @[ICache.scala 225:33]
  wire  s1_tag_hit_3; // @[ICache.scala 225:26]
  wire  _T_146; // @[ICache.scala 140:35]
  reg  s2_valid; // @[ICache.scala 140:25]
  reg [31:0] _RAND_38;
  reg  s2_hit; // @[ICache.scala 141:23]
  reg [31:0] _RAND_39;
  reg  invalidated; // @[ICache.scala 143:24]
  reg [31:0] _RAND_40;
  reg  refill_valid; // @[ICache.scala 144:29]
  reg [31:0] _RAND_41;
  wire  _T_156; // @[ICache.scala 148:26]
  wire  s2_miss; // @[ICache.scala 148:37]
  reg  _T_160; // @[ICache.scala 150:45]
  reg [31:0] _RAND_42;
  wire  s2_request_refill; // @[ICache.scala 150:35]
  wire  refill_fire; // @[Decoupled.scala 37:37]
  wire  _T_158; // @[ICache.scala 149:41]
  wire  s1_can_request_refill; // @[ICache.scala 149:31]
  wire  _T_161; // @[ICache.scala 151:53]
  reg [31:0] refill_addr; // @[Reg.scala 11:16]
  reg [31:0] _RAND_43;
  wire [19:0] refill_tag; // @[ICache.scala 152:31]
  wire [5:0] refill_idx; // @[ICache.scala 153:31]
  wire  refill_one_beat; // @[ICache.scala 154:41]
  wire  s0_valid; // @[Decoupled.scala 37:37]
  wire [26:0] _T_170; // @[package.scala 185:77]
  wire [8:0] _T_173; // @[Edges.scala 220:59]
  wire [8:0] _T_175; // @[Edges.scala 221:14]
  reg [8:0] _T_177; // @[Edges.scala 229:27]
  reg [31:0] _RAND_44;
  wire [8:0] _T_180; // @[Edges.scala 230:28]
  wire  _T_181; // @[Edges.scala 231:25]
  wire  _T_182; // @[Edges.scala 232:25]
  wire  _T_183; // @[Edges.scala 232:47]
  wire  _T_184; // @[Edges.scala 232:37]
  wire  d_done; // @[Edges.scala 233:22]
  wire [8:0] refill_cnt; // @[Edges.scala 234:25]
  wire  refill_done; // @[ICache.scala 162:37]
  reg [15:0] _T_189; // @[LFSR.scala 22:23]
  reg [31:0] _RAND_45;
  wire  _T_192; // @[LFSR.scala 23:43]
  wire  _T_194; // @[LFSR.scala 23:51]
  wire  _T_196; // @[LFSR.scala 23:59]
  wire [15:0] _T_198; // @[Cat.scala 30:58]
  wire [1:0] repl_way; // @[ICache.scala 168:33]
  wire [7:0] _T_201; // @[Cat.scala 30:58]
  wire  _T_271; // @[ICache.scala 198:72]
  wire [255:0] _T_272; // @[ICache.scala 198:32]
  wire [255:0] _T_273; // @[ICache.scala 198:32]
  wire [255:0] _T_275; // @[ICache.scala 198:32]
  wire  _GEN_28; // @[ICache.scala 201:21]
  wire  s1_tl_error_0; // @[ICache.scala 227:32]
  wire  s1_tl_error_1; // @[ICache.scala 227:32]
  wire  s1_tl_error_2; // @[ICache.scala 227:32]
  wire  s1_tl_error_3; // @[ICache.scala 227:32]
  wire [1:0] _T_430; // @[Bitwise.scala 48:55]
  wire [1:0] _T_431; // @[Bitwise.scala 48:55]
  wire [2:0] _T_432; // @[Bitwise.scala 48:55]
  wire  _T_433; // @[ICache.scala 230:115]
  wire  _T_434; // @[ICache.scala 230:39]
  wire  _T_436; // @[ICache.scala 230:9]
  wire  _T_460; // @[ICache.scala 247:28]
  wire  _T_465; // @[ICache.scala 248:32]
  wire [8:0] _T_470; // @[ICache.scala 249:52]
  wire [8:0] _T_471; // @[ICache.scala 249:79]
  wire [31:0] _GEN_52; // @[ICache.scala 259:71]
  wire [31:0] _GEN_53; // @[ICache.scala 259:71]
  wire [31:0] _GEN_54; // @[ICache.scala 259:71]
  wire [31:0] _GEN_55; // @[ICache.scala 259:71]
  wire  _T_530; // @[ICache.scala 247:28]
  reg  s2_tag_hit_0; // @[Reg.scala 11:16]
  reg [31:0] _RAND_46;
  reg  s2_tag_hit_1; // @[Reg.scala 11:16]
  reg [31:0] _RAND_47;
  reg  s2_tag_hit_2; // @[Reg.scala 11:16]
  reg [31:0] _RAND_48;
  reg  s2_tag_hit_3; // @[Reg.scala 11:16]
  reg [31:0] _RAND_49;
  reg [31:0] s2_dout_0; // @[Reg.scala 11:16]
  reg [31:0] _RAND_50;
  reg [31:0] s2_dout_1; // @[Reg.scala 11:16]
  reg [31:0] _RAND_51;
  reg [31:0] s2_dout_2; // @[Reg.scala 11:16]
  reg [31:0] _RAND_52;
  reg [31:0] s2_dout_3; // @[Reg.scala 11:16]
  reg [31:0] _RAND_53;
  wire [31:0] _T_666; // @[Mux.scala 19:72]
  wire [31:0] _T_667; // @[Mux.scala 19:72]
  wire [31:0] _T_668; // @[Mux.scala 19:72]
  wire [31:0] _T_669; // @[Mux.scala 19:72]
  wire [31:0] _T_670; // @[Mux.scala 19:72]
  wire [31:0] _T_671; // @[Mux.scala 19:72]
  wire [3:0] _T_708; // @[ICache.scala 272:43]
  wire  _T_709; // @[ICache.scala 272:50]
  reg  s2_tl_error; // @[Reg.scala 11:16]
  reg [31:0] _RAND_54;
  wire  _GEN_99; // @[ICache.scala 419:22]
  reg [6:0] ICache_state; // @[Register tracking ICache state]
  reg [31:0] _RAND_55;
  reg  ICache_cov [0:127]; // @[Coverage map for ICache]
  reg [31:0] _RAND_56;
  wire  ICache_cov_read_data; // @[Coverage map for ICache]
  wire [6:0] ICache_cov_read_addr; // @[Coverage map for ICache]
  wire  ICache_cov_write_data; // @[Coverage map for ICache]
  wire [6:0] ICache_cov_write_addr; // @[Coverage map for ICache]
  wire  ICache_cov_write_mask; // @[Coverage map for ICache]
  wire  ICache_cov_write_en; // @[Coverage map for ICache]
  reg [29:0] ICache_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_57;
  wire  s2_hit_shl;
  wire [6:0] s2_hit_pad;
  wire [1:0] s2_valid_shl;
  wire [6:0] s2_valid_pad;
  wire [2:0] refill_valid_shl;
  wire [6:0] refill_valid_pad;
  wire [3:0] invalidated_shl;
  wire [6:0] invalidated_pad;
  wire [4:0] _T_160_shl;
  wire [6:0] _T_160_pad;
  wire [5:0] s1_valid_shl;
  wire [6:0] s1_valid_pad;
  wire [6:0] s2_tag_hit_0_shl;
  wire [6:0] s2_tag_hit_0_pad;
  wire [6:0] s2_tag_hit_1_shl;
  wire [6:0] s2_tag_hit_1_pad;
  wire [6:0] s2_tag_hit_2_shl;
  wire [6:0] s2_tag_hit_2_pad;
  wire [6:0] s2_tag_hit_3_shl;
  wire [6:0] s2_tag_hit_3_pad;
  wire [6:0] ICache_xor3;
  wire [6:0] ICache_xor10;
  wire [6:0] ICache_xor4;
  wire [6:0] ICache_xor1;
  wire [6:0] ICache_xor5;
  wire [6:0] ICache_xor14;
  wire [6:0] ICache_xor6;
  wire [6:0] ICache_xor2;
  wire [6:0] ICache_xor0;
  wire  stopEn0;
  reg  ICache_metaAssert;
  reg [31:0] _RAND_58;
  assign tag_array_0_tag_rdata_addr = tag_array_0_tag_rdata_addr_pipe_0;
  assign tag_array_0_tag_rdata_data = tag_array_0[tag_array_0_tag_rdata_addr]; // @[DescribedSRAM.scala 23:21]
  assign tag_array_0__T_256_data = {auto_master_out_d_bits_corrupt,refill_tag};
  assign tag_array_0__T_256_addr = refill_addr[11:6];
  assign tag_array_0__T_256_mask = repl_way == 2'h0;
  assign tag_array_0__T_256_en = refill_one_beat & d_done;
  assign tag_array_1_tag_rdata_addr = tag_array_1_tag_rdata_addr_pipe_0;
  assign tag_array_1_tag_rdata_data = tag_array_1[tag_array_1_tag_rdata_addr]; // @[DescribedSRAM.scala 23:21]
  assign tag_array_1__T_256_data = {auto_master_out_d_bits_corrupt,refill_tag};
  assign tag_array_1__T_256_addr = refill_addr[11:6];
  assign tag_array_1__T_256_mask = repl_way == 2'h1;
  assign tag_array_1__T_256_en = refill_one_beat & d_done;
  assign tag_array_2_tag_rdata_addr = tag_array_2_tag_rdata_addr_pipe_0;
  assign tag_array_2_tag_rdata_data = tag_array_2[tag_array_2_tag_rdata_addr]; // @[DescribedSRAM.scala 23:21]
  assign tag_array_2__T_256_data = {auto_master_out_d_bits_corrupt,refill_tag};
  assign tag_array_2__T_256_addr = refill_addr[11:6];
  assign tag_array_2__T_256_mask = repl_way == 2'h2;
  assign tag_array_2__T_256_en = refill_one_beat & d_done;
  assign tag_array_3_tag_rdata_addr = tag_array_3_tag_rdata_addr_pipe_0;
  assign tag_array_3_tag_rdata_data = tag_array_3[tag_array_3_tag_rdata_addr]; // @[DescribedSRAM.scala 23:21]
  assign tag_array_3__T_256_data = {auto_master_out_d_bits_corrupt,refill_tag};
  assign tag_array_3__T_256_addr = refill_addr[11:6];
  assign tag_array_3__T_256_mask = repl_way == 2'h3;
  assign tag_array_3__T_256_en = refill_one_beat & d_done;
  assign data_arrays_0_0__T_513_addr = data_arrays_0_0__T_513_addr_pipe_0;
  assign data_arrays_0_0__T_513_data = data_arrays_0_0[data_arrays_0_0__T_513_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_0__T_495_data = auto_master_out_d_bits_data[31:0];
  assign data_arrays_0_0__T_495_addr = refill_one_beat ? _T_471 : io_req_bits_addr[11:3];
  assign data_arrays_0_0__T_495_mask = repl_way == 2'h0;
  assign data_arrays_0_0__T_495_en = refill_one_beat & ~invalidated;
  assign data_arrays_0_1__T_513_addr = data_arrays_0_1__T_513_addr_pipe_0;
  assign data_arrays_0_1__T_513_data = data_arrays_0_1[data_arrays_0_1__T_513_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_1__T_495_data = auto_master_out_d_bits_data[31:0];
  assign data_arrays_0_1__T_495_addr = refill_one_beat ? _T_471 : io_req_bits_addr[11:3];
  assign data_arrays_0_1__T_495_mask = repl_way == 2'h1;
  assign data_arrays_0_1__T_495_en = refill_one_beat & ~invalidated;
  assign data_arrays_0_2__T_513_addr = data_arrays_0_2__T_513_addr_pipe_0;
  assign data_arrays_0_2__T_513_data = data_arrays_0_2[data_arrays_0_2__T_513_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_2__T_495_data = auto_master_out_d_bits_data[31:0];
  assign data_arrays_0_2__T_495_addr = refill_one_beat ? _T_471 : io_req_bits_addr[11:3];
  assign data_arrays_0_2__T_495_mask = repl_way == 2'h2;
  assign data_arrays_0_2__T_495_en = refill_one_beat & ~invalidated;
  assign data_arrays_0_3__T_513_addr = data_arrays_0_3__T_513_addr_pipe_0;
  assign data_arrays_0_3__T_513_data = data_arrays_0_3[data_arrays_0_3__T_513_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_0_3__T_495_data = auto_master_out_d_bits_data[31:0];
  assign data_arrays_0_3__T_495_addr = refill_one_beat ? _T_471 : io_req_bits_addr[11:3];
  assign data_arrays_0_3__T_495_mask = repl_way == 2'h3;
  assign data_arrays_0_3__T_495_en = refill_one_beat & ~invalidated;
  assign data_arrays_1_0__T_583_addr = data_arrays_1_0__T_583_addr_pipe_0;
  assign data_arrays_1_0__T_583_data = data_arrays_1_0[data_arrays_1_0__T_583_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_1_0__T_565_data = auto_master_out_d_bits_data[63:32];
  assign data_arrays_1_0__T_565_addr = refill_one_beat ? _T_471 : io_req_bits_addr[11:3];
  assign data_arrays_1_0__T_565_mask = repl_way == 2'h0;
  assign data_arrays_1_0__T_565_en = refill_one_beat & ~invalidated;
  assign data_arrays_1_1__T_583_addr = data_arrays_1_1__T_583_addr_pipe_0;
  assign data_arrays_1_1__T_583_data = data_arrays_1_1[data_arrays_1_1__T_583_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_1_1__T_565_data = auto_master_out_d_bits_data[63:32];
  assign data_arrays_1_1__T_565_addr = refill_one_beat ? _T_471 : io_req_bits_addr[11:3];
  assign data_arrays_1_1__T_565_mask = repl_way == 2'h1;
  assign data_arrays_1_1__T_565_en = refill_one_beat & ~invalidated;
  assign data_arrays_1_2__T_583_addr = data_arrays_1_2__T_583_addr_pipe_0;
  assign data_arrays_1_2__T_583_data = data_arrays_1_2[data_arrays_1_2__T_583_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_1_2__T_565_data = auto_master_out_d_bits_data[63:32];
  assign data_arrays_1_2__T_565_addr = refill_one_beat ? _T_471 : io_req_bits_addr[11:3];
  assign data_arrays_1_2__T_565_mask = repl_way == 2'h2;
  assign data_arrays_1_2__T_565_en = refill_one_beat & ~invalidated;
  assign data_arrays_1_3__T_583_addr = data_arrays_1_3__T_583_addr_pipe_0;
  assign data_arrays_1_3__T_583_data = data_arrays_1_3[data_arrays_1_3__T_583_addr]; // @[DescribedSRAM.scala 23:21]
  assign data_arrays_1_3__T_565_data = auto_master_out_d_bits_data[63:32];
  assign data_arrays_1_3__T_565_addr = refill_one_beat ? _T_471 : io_req_bits_addr[11:3];
  assign data_arrays_1_3__T_565_mask = repl_way == 2'h3;
  assign data_arrays_1_3__T_565_en = refill_one_beat & ~invalidated;
  assign _T_322 = {1'h0,io_s1_paddr[11:6]}; // @[Cat.scala 30:58]
  assign _T_323 = vb_array >> _T_322; // @[ICache.scala 222:25]
  assign _T_329 = tag_array_0_tag_rdata_data[19:0] == io_s1_paddr[31:12]; // @[ICache.scala 225:33]
  assign s1_tag_hit_0 = _T_323[0] & _T_329; // @[ICache.scala 225:26]
  assign _T_350 = {1'h1,io_s1_paddr[11:6]}; // @[Cat.scala 30:58]
  assign _T_351 = vb_array >> _T_350; // @[ICache.scala 222:25]
  assign _T_357 = tag_array_1_tag_rdata_data[19:0] == io_s1_paddr[31:12]; // @[ICache.scala 225:33]
  assign s1_tag_hit_1 = _T_351[0] & _T_357; // @[ICache.scala 225:26]
  assign _T_141 = s1_tag_hit_0 | s1_tag_hit_1; // @[ICache.scala 138:35]
  assign _T_378 = {2'h2,io_s1_paddr[11:6]}; // @[Cat.scala 30:58]
  assign _T_379 = vb_array >> _T_378; // @[ICache.scala 222:25]
  assign _T_385 = tag_array_2_tag_rdata_data[19:0] == io_s1_paddr[31:12]; // @[ICache.scala 225:33]
  assign s1_tag_hit_2 = _T_379[0] & _T_385; // @[ICache.scala 225:26]
  assign _T_142 = _T_141 | s1_tag_hit_2; // @[ICache.scala 138:35]
  assign _T_406 = {2'h3,io_s1_paddr[11:6]}; // @[Cat.scala 30:58]
  assign _T_407 = vb_array >> _T_406; // @[ICache.scala 222:25]
  assign _T_413 = tag_array_3_tag_rdata_data[19:0] == io_s1_paddr[31:12]; // @[ICache.scala 225:33]
  assign s1_tag_hit_3 = _T_407[0] & _T_413; // @[ICache.scala 225:26]
  assign _T_146 = s1_valid & ~io_s1_kill; // @[ICache.scala 140:35]
  assign _T_156 = s2_valid & ~s2_hit; // @[ICache.scala 148:26]
  assign s2_miss = _T_156 & ~io_s2_kill; // @[ICache.scala 148:37]
  assign s2_request_refill = s2_miss & _T_160; // @[ICache.scala 150:35]
  assign refill_fire = auto_master_out_a_ready & s2_request_refill; // @[Decoupled.scala 37:37]
  assign _T_158 = s2_miss | refill_valid; // @[ICache.scala 149:41]
  assign s1_can_request_refill = ~_T_158; // @[ICache.scala 149:31]
  assign _T_161 = s1_valid & s1_can_request_refill; // @[ICache.scala 151:53]
  assign refill_tag = refill_addr[31:12]; // @[ICache.scala 152:31]
  assign refill_idx = refill_addr[11:6]; // @[ICache.scala 153:31]
  assign refill_one_beat = auto_master_out_d_valid & auto_master_out_d_bits_opcode[0]; // @[ICache.scala 154:41]
  assign s0_valid = io_req_ready & io_req_valid; // @[Decoupled.scala 37:37]
  assign _T_170 = 27'hfff << auto_master_out_d_bits_size; // @[package.scala 185:77]
  assign _T_173 = ~_T_170[11:3]; // @[Edges.scala 220:59]
  assign _T_175 = auto_master_out_d_bits_opcode[0] ? _T_173 : 9'h0; // @[Edges.scala 221:14]
  assign _T_180 = _T_177 - 9'h1; // @[Edges.scala 230:28]
  assign _T_181 = _T_177 == 9'h0; // @[Edges.scala 231:25]
  assign _T_182 = _T_177 == 9'h1; // @[Edges.scala 232:25]
  assign _T_183 = _T_175 == 9'h0; // @[Edges.scala 232:47]
  assign _T_184 = _T_182 | _T_183; // @[Edges.scala 232:37]
  assign d_done = _T_184 & auto_master_out_d_valid; // @[Edges.scala 233:22]
  assign refill_cnt = _T_175 & ~_T_180; // @[Edges.scala 234:25]
  assign refill_done = refill_one_beat & d_done; // @[ICache.scala 162:37]
  assign _T_192 = _T_189[0] ^ _T_189[2]; // @[LFSR.scala 23:43]
  assign _T_194 = _T_192 ^ _T_189[3]; // @[LFSR.scala 23:51]
  assign _T_196 = _T_194 ^ _T_189[5]; // @[LFSR.scala 23:59]
  assign _T_198 = {_T_196,_T_189[15:1]}; // @[Cat.scala 30:58]
  assign repl_way = _T_189[1:0]; // @[ICache.scala 168:33]
  assign _T_201 = {repl_way,refill_idx}; // @[Cat.scala 30:58]
  assign _T_271 = refill_done & ~invalidated; // @[ICache.scala 198:72]
  assign _T_272 = 256'h1 << _T_201; // @[ICache.scala 198:32]
  assign _T_273 = vb_array | _T_272; // @[ICache.scala 198:32]
  assign _T_275 = ~vb_array | _T_272; // @[ICache.scala 198:32]
  assign _GEN_28 = io_invalidate | invalidated; // @[ICache.scala 201:21]
  assign s1_tl_error_0 = s1_tag_hit_0 & tag_array_0_tag_rdata_data[20]; // @[ICache.scala 227:32]
  assign s1_tl_error_1 = s1_tag_hit_1 & tag_array_1_tag_rdata_data[20]; // @[ICache.scala 227:32]
  assign s1_tl_error_2 = s1_tag_hit_2 & tag_array_2_tag_rdata_data[20]; // @[ICache.scala 227:32]
  assign s1_tl_error_3 = s1_tag_hit_3 & tag_array_3_tag_rdata_data[20]; // @[ICache.scala 227:32]
  assign _T_430 = s1_tag_hit_0 + s1_tag_hit_1; // @[Bitwise.scala 48:55]
  assign _T_431 = s1_tag_hit_2 + s1_tag_hit_3; // @[Bitwise.scala 48:55]
  assign _T_432 = _T_430 + _T_431; // @[Bitwise.scala 48:55]
  assign _T_433 = _T_432 <= 3'h1; // @[ICache.scala 230:115]
  assign _T_434 = ~s1_valid | _T_433; // @[ICache.scala 230:39]
  assign _T_436 = _T_434 | reset; // @[ICache.scala 230:9]
  assign _T_460 = s0_valid & ~io_req_bits_addr[2]; // @[ICache.scala 247:28]
  assign _T_465 = refill_one_beat & ~invalidated; // @[ICache.scala 248:32]
  assign _T_470 = {refill_idx, 3'h0}; // @[ICache.scala 249:52]
  assign _T_471 = _T_470 | refill_cnt; // @[ICache.scala 249:79]
  assign _GEN_52 = data_arrays_0_0__T_513_data; // @[ICache.scala 259:71]
  assign _GEN_53 = data_arrays_0_1__T_513_data; // @[ICache.scala 259:71]
  assign _GEN_54 = data_arrays_0_2__T_513_data; // @[ICache.scala 259:71]
  assign _GEN_55 = data_arrays_0_3__T_513_data; // @[ICache.scala 259:71]
  assign _T_530 = s0_valid & io_req_bits_addr[2]; // @[ICache.scala 247:28]
  assign _T_666 = s2_tag_hit_0 ? s2_dout_0 : 32'h0; // @[Mux.scala 19:72]
  assign _T_667 = s2_tag_hit_1 ? s2_dout_1 : 32'h0; // @[Mux.scala 19:72]
  assign _T_668 = s2_tag_hit_2 ? s2_dout_2 : 32'h0; // @[Mux.scala 19:72]
  assign _T_669 = s2_tag_hit_3 ? s2_dout_3 : 32'h0; // @[Mux.scala 19:72]
  assign _T_670 = _T_666 | _T_667; // @[Mux.scala 19:72]
  assign _T_671 = _T_670 | _T_668; // @[Mux.scala 19:72]
  assign _T_708 = {s1_tl_error_3,s1_tl_error_2,s1_tl_error_1,s1_tl_error_0}; // @[ICache.scala 272:43]
  assign _T_709 = _T_708 != 4'h0; // @[ICache.scala 272:50]
  assign _GEN_99 = refill_fire | refill_valid; // @[ICache.scala 419:22]
  assign auto_master_out_a_valid = s2_miss & _T_160; // @[LazyModule.scala 173:49]
  assign auto_master_out_a_bits_address = {refill_addr[31:6], 6'h0}; // @[LazyModule.scala 173:49]
  assign io_req_ready = ~refill_one_beat; // @[ICache.scala 156:16]
  assign io_resp_valid = s2_valid & s2_hit; // @[ICache.scala 299:21]
  assign io_resp_bits_data = _T_671 | _T_669; // @[ICache.scala 296:25]
  assign io_resp_bits_ae = s2_tl_error; // @[ICache.scala 297:23]
  assign ICache_cov_read_addr = ICache_state;
  assign ICache_cov_read_data = ICache_cov[ICache_cov_read_addr]; // @[Coverage map for ICache]
  assign ICache_cov_write_data = 1'h1;
  assign ICache_cov_write_addr = ICache_state;
  assign ICache_cov_write_mask = 1'h1;
  assign ICache_cov_write_en = 1'h1;
  assign s2_hit_shl = s2_hit;
  assign s2_hit_pad = {6'h0,s2_hit_shl};
  assign s2_valid_shl = {s2_valid, 1'h0};
  assign s2_valid_pad = {5'h0,s2_valid_shl};
  assign refill_valid_shl = {refill_valid, 2'h0};
  assign refill_valid_pad = {4'h0,refill_valid_shl};
  assign invalidated_shl = {invalidated, 3'h0};
  assign invalidated_pad = {3'h0,invalidated_shl};
  assign _T_160_shl = {_T_160, 4'h0};
  assign _T_160_pad = {2'h0,_T_160_shl};
  assign s1_valid_shl = {s1_valid, 5'h0};
  assign s1_valid_pad = {1'h0,s1_valid_shl};
  assign s2_tag_hit_0_shl = {s2_tag_hit_0, 6'h0};
  assign s2_tag_hit_0_pad = s2_tag_hit_0_shl;
  assign s2_tag_hit_1_shl = {s2_tag_hit_1, 6'h0};
  assign s2_tag_hit_1_pad = s2_tag_hit_1_shl;
  assign s2_tag_hit_2_shl = {s2_tag_hit_2, 6'h0};
  assign s2_tag_hit_2_pad = s2_tag_hit_2_shl;
  assign s2_tag_hit_3_shl = {s2_tag_hit_3, 6'h0};
  assign s2_tag_hit_3_pad = s2_tag_hit_3_shl;
  assign ICache_xor3 = s2_hit_pad ^ s2_valid_pad;
  assign ICache_xor10 = invalidated_pad ^ _T_160_pad;
  assign ICache_xor4 = refill_valid_pad ^ ICache_xor10;
  assign ICache_xor1 = ICache_xor3 ^ ICache_xor4;
  assign ICache_xor5 = s1_valid_pad ^ s2_tag_hit_0_pad;
  assign ICache_xor14 = s2_tag_hit_2_pad ^ s2_tag_hit_3_pad;
  assign ICache_xor6 = s2_tag_hit_1_pad ^ ICache_xor14;
  assign ICache_xor2 = ICache_xor5 ^ ICache_xor6;
  assign ICache_xor0 = ICache_xor1 ^ ICache_xor2;
  assign io_covSum = ICache_covSum;
  assign stopEn0 = ~_T_436;
  assign metaAssert = ICache_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_0[initvar] = _RAND_0[20:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tag_array_0_tag_rdata_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  tag_array_0_tag_rdata_addr_pipe_0 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_1[initvar] = _RAND_3[20:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  tag_array_1_tag_rdata_en_pipe_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  tag_array_1_tag_rdata_addr_pipe_0 = _RAND_5[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_2[initvar] = _RAND_6[20:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  tag_array_2_tag_rdata_en_pipe_0 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  tag_array_2_tag_rdata_addr_pipe_0 = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_3[initvar] = _RAND_9[20:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  tag_array_3_tag_rdata_en_pipe_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  tag_array_3_tag_rdata_addr_pipe_0 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_0[initvar] = _RAND_12[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  data_arrays_0_0__T_513_en_pipe_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  data_arrays_0_0__T_513_addr_pipe_0 = _RAND_14[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_1[initvar] = _RAND_15[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  data_arrays_0_1__T_513_en_pipe_0 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  data_arrays_0_1__T_513_addr_pipe_0 = _RAND_17[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_2[initvar] = _RAND_18[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  data_arrays_0_2__T_513_en_pipe_0 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  data_arrays_0_2__T_513_addr_pipe_0 = _RAND_20[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_3[initvar] = _RAND_21[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  data_arrays_0_3__T_513_en_pipe_0 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  data_arrays_0_3__T_513_addr_pipe_0 = _RAND_23[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_1_0[initvar] = _RAND_24[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  data_arrays_1_0__T_583_en_pipe_0 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  data_arrays_1_0__T_583_addr_pipe_0 = _RAND_26[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_1_1[initvar] = _RAND_27[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  data_arrays_1_1__T_583_en_pipe_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  data_arrays_1_1__T_583_addr_pipe_0 = _RAND_29[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_1_2[initvar] = _RAND_30[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  data_arrays_1_2__T_583_en_pipe_0 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  data_arrays_1_2__T_583_addr_pipe_0 = _RAND_32[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_1_3[initvar] = _RAND_33[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  data_arrays_1_3__T_583_en_pipe_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  data_arrays_1_3__T_583_addr_pipe_0 = _RAND_35[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  s1_valid = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {8{`RANDOM}};
  vb_array = _RAND_37[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  s2_valid = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  s2_hit = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  invalidated = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  refill_valid = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_160 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  refill_addr = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_177 = _RAND_44[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_189 = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  s2_tag_hit_0 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  s2_tag_hit_1 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  s2_tag_hit_2 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  s2_tag_hit_3 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  s2_dout_0 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  s2_dout_1 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  s2_dout_2 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  s2_dout_3 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  s2_tl_error = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  ICache_state = _RAND_55[6:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ICache_cov[initvar] = _RAND_56[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  ICache_covSum = _RAND_57[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  ICache_metaAssert = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(tag_array_0__T_256_en & tag_array_0__T_256_mask) begin
      tag_array_0[tag_array_0__T_256_addr] <= tag_array_0__T_256_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      tag_array_0_tag_rdata_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_0_tag_rdata_en_pipe_0 <= ~refill_done & s0_valid;
    end
    if (metaReset) begin
      tag_array_0_tag_rdata_addr_pipe_0 <= 6'h0;
    end else if (~refill_done & s0_valid) begin
      tag_array_0_tag_rdata_addr_pipe_0 <= io_req_bits_addr[11:6];
    end
    if(tag_array_1__T_256_en & tag_array_1__T_256_mask) begin
      tag_array_1[tag_array_1__T_256_addr] <= tag_array_1__T_256_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      tag_array_1_tag_rdata_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_1_tag_rdata_en_pipe_0 <= ~refill_done & s0_valid;
    end
    if (metaReset) begin
      tag_array_1_tag_rdata_addr_pipe_0 <= 6'h0;
    end else if (~refill_done & s0_valid) begin
      tag_array_1_tag_rdata_addr_pipe_0 <= io_req_bits_addr[11:6];
    end
    if(tag_array_2__T_256_en & tag_array_2__T_256_mask) begin
      tag_array_2[tag_array_2__T_256_addr] <= tag_array_2__T_256_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      tag_array_2_tag_rdata_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_2_tag_rdata_en_pipe_0 <= ~refill_done & s0_valid;
    end
    if (metaReset) begin
      tag_array_2_tag_rdata_addr_pipe_0 <= 6'h0;
    end else if (~refill_done & s0_valid) begin
      tag_array_2_tag_rdata_addr_pipe_0 <= io_req_bits_addr[11:6];
    end
    if(tag_array_3__T_256_en & tag_array_3__T_256_mask) begin
      tag_array_3[tag_array_3__T_256_addr] <= tag_array_3__T_256_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      tag_array_3_tag_rdata_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_3_tag_rdata_en_pipe_0 <= ~refill_done & s0_valid;
    end
    if (metaReset) begin
      tag_array_3_tag_rdata_addr_pipe_0 <= 6'h0;
    end else if (~refill_done & s0_valid) begin
      tag_array_3_tag_rdata_addr_pipe_0 <= io_req_bits_addr[11:6];
    end
    if(data_arrays_0_0__T_495_en & data_arrays_0_0__T_495_mask) begin
      data_arrays_0_0[data_arrays_0_0__T_495_addr] <= data_arrays_0_0__T_495_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_0__T_513_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_0__T_513_en_pipe_0 <= ~_T_465 & _T_460;
    end
    if (metaReset) begin
      data_arrays_0_0__T_513_addr_pipe_0 <= 9'h0;
    end else if (~_T_465 & _T_460) begin
      if (refill_one_beat) begin
        data_arrays_0_0__T_513_addr_pipe_0 <= _T_471;
      end else begin
        data_arrays_0_0__T_513_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if(data_arrays_0_1__T_495_en & data_arrays_0_1__T_495_mask) begin
      data_arrays_0_1[data_arrays_0_1__T_495_addr] <= data_arrays_0_1__T_495_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_1__T_513_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_1__T_513_en_pipe_0 <= ~_T_465 & _T_460;
    end
    if (metaReset) begin
      data_arrays_0_1__T_513_addr_pipe_0 <= 9'h0;
    end else if (~_T_465 & _T_460) begin
      if (refill_one_beat) begin
        data_arrays_0_1__T_513_addr_pipe_0 <= _T_471;
      end else begin
        data_arrays_0_1__T_513_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if(data_arrays_0_2__T_495_en & data_arrays_0_2__T_495_mask) begin
      data_arrays_0_2[data_arrays_0_2__T_495_addr] <= data_arrays_0_2__T_495_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_2__T_513_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_2__T_513_en_pipe_0 <= ~_T_465 & _T_460;
    end
    if (metaReset) begin
      data_arrays_0_2__T_513_addr_pipe_0 <= 9'h0;
    end else if (~_T_465 & _T_460) begin
      if (refill_one_beat) begin
        data_arrays_0_2__T_513_addr_pipe_0 <= _T_471;
      end else begin
        data_arrays_0_2__T_513_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if(data_arrays_0_3__T_495_en & data_arrays_0_3__T_495_mask) begin
      data_arrays_0_3[data_arrays_0_3__T_495_addr] <= data_arrays_0_3__T_495_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_0_3__T_513_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_3__T_513_en_pipe_0 <= ~_T_465 & _T_460;
    end
    if (metaReset) begin
      data_arrays_0_3__T_513_addr_pipe_0 <= 9'h0;
    end else if (~_T_465 & _T_460) begin
      if (refill_one_beat) begin
        data_arrays_0_3__T_513_addr_pipe_0 <= _T_471;
      end else begin
        data_arrays_0_3__T_513_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if(data_arrays_1_0__T_565_en & data_arrays_1_0__T_565_mask) begin
      data_arrays_1_0[data_arrays_1_0__T_565_addr] <= data_arrays_1_0__T_565_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_1_0__T_583_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_1_0__T_583_en_pipe_0 <= ~_T_465 & _T_530;
    end
    if (metaReset) begin
      data_arrays_1_0__T_583_addr_pipe_0 <= 9'h0;
    end else if (~_T_465 & _T_530) begin
      if (refill_one_beat) begin
        data_arrays_1_0__T_583_addr_pipe_0 <= _T_471;
      end else begin
        data_arrays_1_0__T_583_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if(data_arrays_1_1__T_565_en & data_arrays_1_1__T_565_mask) begin
      data_arrays_1_1[data_arrays_1_1__T_565_addr] <= data_arrays_1_1__T_565_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_1_1__T_583_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_1_1__T_583_en_pipe_0 <= ~_T_465 & _T_530;
    end
    if (metaReset) begin
      data_arrays_1_1__T_583_addr_pipe_0 <= 9'h0;
    end else if (~_T_465 & _T_530) begin
      if (refill_one_beat) begin
        data_arrays_1_1__T_583_addr_pipe_0 <= _T_471;
      end else begin
        data_arrays_1_1__T_583_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if(data_arrays_1_2__T_565_en & data_arrays_1_2__T_565_mask) begin
      data_arrays_1_2[data_arrays_1_2__T_565_addr] <= data_arrays_1_2__T_565_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_1_2__T_583_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_1_2__T_583_en_pipe_0 <= ~_T_465 & _T_530;
    end
    if (metaReset) begin
      data_arrays_1_2__T_583_addr_pipe_0 <= 9'h0;
    end else if (~_T_465 & _T_530) begin
      if (refill_one_beat) begin
        data_arrays_1_2__T_583_addr_pipe_0 <= _T_471;
      end else begin
        data_arrays_1_2__T_583_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if(data_arrays_1_3__T_565_en & data_arrays_1_3__T_565_mask) begin
      data_arrays_1_3[data_arrays_1_3__T_565_addr] <= data_arrays_1_3__T_565_data; // @[DescribedSRAM.scala 23:21]
    end
    if (metaReset) begin
      data_arrays_1_3__T_583_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_1_3__T_583_en_pipe_0 <= ~_T_465 & _T_530;
    end
    if (metaReset) begin
      data_arrays_1_3__T_583_addr_pipe_0 <= 9'h0;
    end else if (~_T_465 & _T_530) begin
      if (refill_one_beat) begin
        data_arrays_1_3__T_583_addr_pipe_0 <= _T_471;
      end else begin
        data_arrays_1_3__T_583_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if (metaReset) begin
      s1_valid <= 1'h0;
    end else if (reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= s0_valid;
    end
    if (metaReset) begin
      vb_array <= 256'h0;
    end else if (reset) begin
      vb_array <= 256'h0;
    end else if (io_invalidate) begin
      vb_array <= 256'h0;
    end else if (refill_one_beat) begin
      if (_T_271) begin
        vb_array <= _T_273;
      end else begin
        vb_array <= ~_T_275;
      end
    end
    if (metaReset) begin
      s2_valid <= 1'h0;
    end else if (reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= _T_146;
    end
    if (metaReset) begin
      s2_hit <= 1'h0;
    end else begin
      s2_hit <= _T_142 | s1_tag_hit_3;
    end
    if (metaReset) begin
      invalidated <= 1'h0;
    end else if (~refill_valid) begin
      invalidated <= 1'h0;
    end else begin
      invalidated <= _GEN_28;
    end
    if (metaReset) begin
      refill_valid <= 1'h0;
    end else if (reset) begin
      refill_valid <= 1'h0;
    end else if (refill_done) begin
      refill_valid <= 1'h0;
    end else begin
      refill_valid <= _GEN_99;
    end
    if (metaReset) begin
      _T_160 <= 1'h0;
    end else begin
      _T_160 <= ~_T_158;
    end
    if (metaReset) begin
      refill_addr <= 32'h0;
    end else if (_T_161) begin
      refill_addr <= io_s1_paddr;
    end
    if (metaReset) begin
      _T_177 <= 9'h0;
    end else if (reset) begin
      _T_177 <= 9'h0;
    end else if (auto_master_out_d_valid) begin
      if (_T_181) begin
        if (auto_master_out_d_bits_opcode[0]) begin
          _T_177 <= _T_173;
        end else begin
          _T_177 <= 9'h0;
        end
      end else begin
        _T_177 <= _T_180;
      end
    end
    if (metaReset) begin
      _T_189 <= 16'h0;
    end else if (reset) begin
      _T_189 <= 16'h1;
    end else if (refill_fire) begin
      _T_189 <= _T_198;
    end
    if (metaReset) begin
      s2_tag_hit_0 <= 1'h0;
    end else if (s1_valid) begin
      s2_tag_hit_0 <= s1_tag_hit_0;
    end
    if (metaReset) begin
      s2_tag_hit_1 <= 1'h0;
    end else if (s1_valid) begin
      s2_tag_hit_1 <= s1_tag_hit_1;
    end
    if (metaReset) begin
      s2_tag_hit_2 <= 1'h0;
    end else if (s1_valid) begin
      s2_tag_hit_2 <= s1_tag_hit_2;
    end
    if (metaReset) begin
      s2_tag_hit_3 <= 1'h0;
    end else if (s1_valid) begin
      s2_tag_hit_3 <= s1_tag_hit_3;
    end
    if (metaReset) begin
      s2_dout_0 <= 32'h0;
    end else if (s1_valid) begin
      if (io_s1_paddr[2]) begin
        s2_dout_0 <= data_arrays_1_0__T_583_data;
      end else begin
        s2_dout_0 <= _GEN_52;
      end
    end
    if (metaReset) begin
      s2_dout_1 <= 32'h0;
    end else if (s1_valid) begin
      if (io_s1_paddr[2]) begin
        s2_dout_1 <= data_arrays_1_1__T_583_data;
      end else begin
        s2_dout_1 <= _GEN_53;
      end
    end
    if (metaReset) begin
      s2_dout_2 <= 32'h0;
    end else if (s1_valid) begin
      if (io_s1_paddr[2]) begin
        s2_dout_2 <= data_arrays_1_2__T_583_data;
      end else begin
        s2_dout_2 <= _GEN_54;
      end
    end
    if (metaReset) begin
      s2_dout_3 <= 32'h0;
    end else if (s1_valid) begin
      if (io_s1_paddr[2]) begin
        s2_dout_3 <= data_arrays_1_3__T_583_data;
      end else begin
        s2_dout_3 <= _GEN_55;
      end
    end
    if (metaReset) begin
      s2_tl_error <= 1'h0;
    end else if (s1_valid) begin
      s2_tl_error <= _T_709;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_436) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ICache.scala:230 assert(!(s1_valid || s1_slaveValid) || PopCount(s1_tag_hit zip s1_tag_disparity map { case (h, d) => h && !d }) <= 1)\n"); // @[ICache.scala 230:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_436) begin
          $fatal; // @[ICache.scala 230:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    ICache_state <= ICache_xor0;
    if (!(ICache_cov_read_data)) begin
      ICache_covSum <= ICache_covSum + 1'h1;
    end
    if (metaReset) begin
      ICache_metaAssert <= 1'h0;
    end else begin
      ICache_metaAssert <= ICache_metaAssert | stopEn0;
    end
  end
  always @(posedge clock) begin
    if(ICache_cov_write_en & ICache_cov_write_mask) begin
      ICache_cov[ICache_cov_write_addr] <= ICache_cov_write_data; // @[Coverage map for ICache]
    end
  end
endmodule
module ShiftQueue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_btb_taken,
  input         io_enq_bits_btb_bridx,
  input  [4:0]  io_enq_bits_btb_entry,
  input  [7:0]  io_enq_bits_btb_bht_history,
  input  [39:0] io_enq_bits_pc,
  input  [31:0] io_enq_bits_data,
  input  [1:0]  io_enq_bits_mask,
  input         io_enq_bits_xcpt_pf_inst,
  input         io_enq_bits_xcpt_ae_inst,
  input         io_enq_bits_replay,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_btb_taken,
  output        io_deq_bits_btb_bridx,
  output [4:0]  io_deq_bits_btb_entry,
  output [7:0]  io_deq_bits_btb_bht_history,
  output [39:0] io_deq_bits_pc,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_xcpt_pf_inst,
  output        io_deq_bits_xcpt_ae_inst,
  output        io_deq_bits_replay,
  output [4:0]  io_mask,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg  _T_60_0; // @[ShiftQueue.scala 20:30]
  reg [31:0] _RAND_0;
  reg  _T_60_1; // @[ShiftQueue.scala 20:30]
  reg [31:0] _RAND_1;
  reg  _T_60_2; // @[ShiftQueue.scala 20:30]
  reg [31:0] _RAND_2;
  reg  _T_60_3; // @[ShiftQueue.scala 20:30]
  reg [31:0] _RAND_3;
  reg  _T_60_4; // @[ShiftQueue.scala 20:30]
  reg [31:0] _RAND_4;
  reg  _T_82_0_btb_taken; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_5;
  reg  _T_82_0_btb_bridx; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_6;
  reg [4:0] _T_82_0_btb_entry; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_7;
  reg [7:0] _T_82_0_btb_bht_history; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_8;
  reg [39:0] _T_82_0_pc; // @[ShiftQueue.scala 21:25]
  reg [63:0] _RAND_9;
  reg [31:0] _T_82_0_data; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_10;
  reg  _T_82_0_xcpt_pf_inst; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_11;
  reg  _T_82_0_xcpt_ae_inst; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_12;
  reg  _T_82_0_replay; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_13;
  reg  _T_82_1_btb_taken; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_14;
  reg  _T_82_1_btb_bridx; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_15;
  reg [4:0] _T_82_1_btb_entry; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_16;
  reg [7:0] _T_82_1_btb_bht_history; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_17;
  reg [39:0] _T_82_1_pc; // @[ShiftQueue.scala 21:25]
  reg [63:0] _RAND_18;
  reg [31:0] _T_82_1_data; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_19;
  reg  _T_82_1_xcpt_pf_inst; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_20;
  reg  _T_82_1_xcpt_ae_inst; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_21;
  reg  _T_82_1_replay; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_22;
  reg  _T_82_2_btb_taken; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_23;
  reg  _T_82_2_btb_bridx; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_24;
  reg [4:0] _T_82_2_btb_entry; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_25;
  reg [7:0] _T_82_2_btb_bht_history; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_26;
  reg [39:0] _T_82_2_pc; // @[ShiftQueue.scala 21:25]
  reg [63:0] _RAND_27;
  reg [31:0] _T_82_2_data; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_28;
  reg  _T_82_2_xcpt_pf_inst; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_29;
  reg  _T_82_2_xcpt_ae_inst; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_30;
  reg  _T_82_2_replay; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_31;
  reg  _T_82_3_btb_taken; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_32;
  reg  _T_82_3_btb_bridx; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_33;
  reg [4:0] _T_82_3_btb_entry; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_34;
  reg [7:0] _T_82_3_btb_bht_history; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_35;
  reg [39:0] _T_82_3_pc; // @[ShiftQueue.scala 21:25]
  reg [63:0] _RAND_36;
  reg [31:0] _T_82_3_data; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_37;
  reg  _T_82_3_xcpt_pf_inst; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_38;
  reg  _T_82_3_xcpt_ae_inst; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_39;
  reg  _T_82_3_replay; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_40;
  reg  _T_82_4_btb_taken; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_41;
  reg  _T_82_4_btb_bridx; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_42;
  reg [4:0] _T_82_4_btb_entry; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_43;
  reg [7:0] _T_82_4_btb_bht_history; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_44;
  reg [39:0] _T_82_4_pc; // @[ShiftQueue.scala 21:25]
  reg [63:0] _RAND_45;
  reg [31:0] _T_82_4_data; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_46;
  reg  _T_82_4_xcpt_pf_inst; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_47;
  reg  _T_82_4_xcpt_ae_inst; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_48;
  reg  _T_82_4_replay; // @[ShiftQueue.scala 21:25]
  reg [31:0] _RAND_49;
  wire  _T_91; // @[Decoupled.scala 37:37]
  wire  _T_93; // @[ShiftQueue.scala 29:45]
  wire  _T_94; // @[ShiftQueue.scala 29:28]
  wire  _T_98; // @[ShiftQueue.scala 30:45]
  wire  _T_99; // @[ShiftQueue.scala 28:10]
  wire  _T_106; // @[ShiftQueue.scala 36:45]
  wire  _T_111; // @[ShiftQueue.scala 29:45]
  wire  _T_112; // @[ShiftQueue.scala 29:28]
  wire  _T_116; // @[ShiftQueue.scala 30:45]
  wire  _T_117; // @[ShiftQueue.scala 28:10]
  wire  _T_124; // @[ShiftQueue.scala 36:45]
  wire  _T_129; // @[ShiftQueue.scala 29:45]
  wire  _T_130; // @[ShiftQueue.scala 29:28]
  wire  _T_134; // @[ShiftQueue.scala 30:45]
  wire  _T_135; // @[ShiftQueue.scala 28:10]
  wire  _T_142; // @[ShiftQueue.scala 36:45]
  wire  _T_147; // @[ShiftQueue.scala 29:45]
  wire  _T_148; // @[ShiftQueue.scala 29:28]
  wire  _T_152; // @[ShiftQueue.scala 30:45]
  wire  _T_153; // @[ShiftQueue.scala 28:10]
  wire  _T_160; // @[ShiftQueue.scala 36:45]
  wire  _T_164; // @[ShiftQueue.scala 29:45]
  wire  _T_169; // @[ShiftQueue.scala 30:45]
  wire  _T_170; // @[ShiftQueue.scala 28:10]
  wire  _T_177; // @[ShiftQueue.scala 36:45]
  wire [1:0] _T_181; // @[ShiftQueue.scala 52:20]
  wire [2:0] _T_183; // @[ShiftQueue.scala 52:20]
  reg  ShiftQueue_state; // @[Register tracking ShiftQueue state]
  reg [31:0] _RAND_50;
  reg  ShiftQueue_cov [0:1]; // @[Coverage map for ShiftQueue]
  reg [31:0] _RAND_51;
  wire  ShiftQueue_cov_read_data; // @[Coverage map for ShiftQueue]
  wire  ShiftQueue_cov_read_addr; // @[Coverage map for ShiftQueue]
  wire  ShiftQueue_cov_write_data; // @[Coverage map for ShiftQueue]
  wire  ShiftQueue_cov_write_addr; // @[Coverage map for ShiftQueue]
  wire  ShiftQueue_cov_write_mask; // @[Coverage map for ShiftQueue]
  wire  ShiftQueue_cov_write_en; // @[Coverage map for ShiftQueue]
  reg [29:0] ShiftQueue_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_52;
  wire  _T_60_3_shl;
  wire  _T_60_3_pad;
  wire  _T_60_0_shl;
  wire  _T_60_0_pad;
  wire  _T_60_4_shl;
  wire  _T_60_4_pad;
  wire  _T_60_1_shl;
  wire  _T_60_1_pad;
  wire  _T_60_2_shl;
  wire  _T_60_2_pad;
  wire  ShiftQueue_xor1;
  wire  ShiftQueue_xor6;
  wire  ShiftQueue_xor2;
  wire  ShiftQueue_xor0;
  assign _T_91 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37]
  assign _T_93 = _T_91 & _T_60_0; // @[ShiftQueue.scala 29:45]
  assign _T_94 = _T_60_1 | _T_93; // @[ShiftQueue.scala 29:28]
  assign _T_98 = _T_91 & ~_T_60_0; // @[ShiftQueue.scala 30:45]
  assign _T_99 = io_deq_ready ? _T_94 : _T_98; // @[ShiftQueue.scala 28:10]
  assign _T_106 = _T_91 | _T_60_0; // @[ShiftQueue.scala 36:45]
  assign _T_111 = _T_91 & _T_60_1; // @[ShiftQueue.scala 29:45]
  assign _T_112 = _T_60_2 | _T_111; // @[ShiftQueue.scala 29:28]
  assign _T_116 = _T_93 & ~_T_60_1; // @[ShiftQueue.scala 30:45]
  assign _T_117 = io_deq_ready ? _T_112 : _T_116; // @[ShiftQueue.scala 28:10]
  assign _T_124 = _T_93 | _T_60_1; // @[ShiftQueue.scala 36:45]
  assign _T_129 = _T_91 & _T_60_2; // @[ShiftQueue.scala 29:45]
  assign _T_130 = _T_60_3 | _T_129; // @[ShiftQueue.scala 29:28]
  assign _T_134 = _T_111 & ~_T_60_2; // @[ShiftQueue.scala 30:45]
  assign _T_135 = io_deq_ready ? _T_130 : _T_134; // @[ShiftQueue.scala 28:10]
  assign _T_142 = _T_111 | _T_60_2; // @[ShiftQueue.scala 36:45]
  assign _T_147 = _T_91 & _T_60_3; // @[ShiftQueue.scala 29:45]
  assign _T_148 = _T_60_4 | _T_147; // @[ShiftQueue.scala 29:28]
  assign _T_152 = _T_129 & ~_T_60_3; // @[ShiftQueue.scala 30:45]
  assign _T_153 = io_deq_ready ? _T_148 : _T_152; // @[ShiftQueue.scala 28:10]
  assign _T_160 = _T_129 | _T_60_3; // @[ShiftQueue.scala 36:45]
  assign _T_164 = _T_91 & _T_60_4; // @[ShiftQueue.scala 29:45]
  assign _T_169 = _T_147 & ~_T_60_4; // @[ShiftQueue.scala 30:45]
  assign _T_170 = io_deq_ready ? _T_164 : _T_169; // @[ShiftQueue.scala 28:10]
  assign _T_177 = _T_147 | _T_60_4; // @[ShiftQueue.scala 36:45]
  assign _T_181 = {_T_60_1,_T_60_0}; // @[ShiftQueue.scala 52:20]
  assign _T_183 = {_T_60_4,_T_60_3,_T_60_2}; // @[ShiftQueue.scala 52:20]
  assign io_enq_ready = ~_T_60_4; // @[ShiftQueue.scala 39:16]
  assign io_deq_valid = io_enq_valid | _T_60_0; // @[ShiftQueue.scala 40:16 ShiftQueue.scala 44:40]
  assign io_deq_bits_btb_taken = _T_60_0 ? _T_82_0_btb_taken : io_enq_bits_btb_taken; // @[ShiftQueue.scala 41:15 ShiftQueue.scala 45:36]
  assign io_deq_bits_btb_bridx = _T_60_0 ? _T_82_0_btb_bridx : io_enq_bits_btb_bridx; // @[ShiftQueue.scala 41:15 ShiftQueue.scala 45:36]
  assign io_deq_bits_btb_entry = _T_60_0 ? _T_82_0_btb_entry : io_enq_bits_btb_entry; // @[ShiftQueue.scala 41:15 ShiftQueue.scala 45:36]
  assign io_deq_bits_btb_bht_history = _T_60_0 ? _T_82_0_btb_bht_history : io_enq_bits_btb_bht_history; // @[ShiftQueue.scala 41:15 ShiftQueue.scala 45:36]
  assign io_deq_bits_pc = _T_60_0 ? _T_82_0_pc : io_enq_bits_pc; // @[ShiftQueue.scala 41:15 ShiftQueue.scala 45:36]
  assign io_deq_bits_data = _T_60_0 ? _T_82_0_data : io_enq_bits_data; // @[ShiftQueue.scala 41:15 ShiftQueue.scala 45:36]
  assign io_deq_bits_xcpt_pf_inst = _T_60_0 ? _T_82_0_xcpt_pf_inst : io_enq_bits_xcpt_pf_inst; // @[ShiftQueue.scala 41:15 ShiftQueue.scala 45:36]
  assign io_deq_bits_xcpt_ae_inst = _T_60_0 ? _T_82_0_xcpt_ae_inst : io_enq_bits_xcpt_ae_inst; // @[ShiftQueue.scala 41:15 ShiftQueue.scala 45:36]
  assign io_deq_bits_replay = _T_60_0 ? _T_82_0_replay : io_enq_bits_replay; // @[ShiftQueue.scala 41:15 ShiftQueue.scala 45:36]
  assign io_mask = {_T_183,_T_181}; // @[ShiftQueue.scala 52:11]
  assign ShiftQueue_cov_read_addr = ShiftQueue_state;
  assign ShiftQueue_cov_read_data = ShiftQueue_cov[ShiftQueue_cov_read_addr]; // @[Coverage map for ShiftQueue]
  assign ShiftQueue_cov_write_data = 1'h1;
  assign ShiftQueue_cov_write_addr = ShiftQueue_state;
  assign ShiftQueue_cov_write_mask = 1'h1;
  assign ShiftQueue_cov_write_en = 1'h1;
  assign _T_60_3_shl = _T_60_3;
  assign _T_60_3_pad = _T_60_3_shl;
  assign _T_60_0_shl = _T_60_0;
  assign _T_60_0_pad = _T_60_0_shl;
  assign _T_60_4_shl = _T_60_4;
  assign _T_60_4_pad = _T_60_4_shl;
  assign _T_60_1_shl = _T_60_1;
  assign _T_60_1_pad = _T_60_1_shl;
  assign _T_60_2_shl = _T_60_2;
  assign _T_60_2_pad = _T_60_2_shl;
  assign ShiftQueue_xor1 = _T_60_3_pad ^ _T_60_0_pad;
  assign ShiftQueue_xor6 = _T_60_1_pad ^ _T_60_2_pad;
  assign ShiftQueue_xor2 = _T_60_4_pad ^ ShiftQueue_xor6;
  assign ShiftQueue_xor0 = ShiftQueue_xor1 ^ ShiftQueue_xor2;
  assign io_covSum = ShiftQueue_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_60_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_60_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_60_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_60_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_60_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_82_0_btb_taken = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_82_0_btb_bridx = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_82_0_btb_entry = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_82_0_btb_bht_history = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {2{`RANDOM}};
  _T_82_0_pc = _RAND_9[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_82_0_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_82_0_xcpt_pf_inst = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_82_0_xcpt_ae_inst = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_82_0_replay = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_82_1_btb_taken = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_82_1_btb_bridx = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_82_1_btb_entry = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_82_1_btb_bht_history = _RAND_17[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {2{`RANDOM}};
  _T_82_1_pc = _RAND_18[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_82_1_data = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_82_1_xcpt_pf_inst = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_82_1_xcpt_ae_inst = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_82_1_replay = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_82_2_btb_taken = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_82_2_btb_bridx = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_82_2_btb_entry = _RAND_25[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_82_2_btb_bht_history = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {2{`RANDOM}};
  _T_82_2_pc = _RAND_27[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_82_2_data = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_82_2_xcpt_pf_inst = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_82_2_xcpt_ae_inst = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_82_2_replay = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_82_3_btb_taken = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_82_3_btb_bridx = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_82_3_btb_entry = _RAND_34[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_82_3_btb_bht_history = _RAND_35[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {2{`RANDOM}};
  _T_82_3_pc = _RAND_36[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_82_3_data = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_82_3_xcpt_pf_inst = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_82_3_xcpt_ae_inst = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_82_3_replay = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_82_4_btb_taken = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_82_4_btb_bridx = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_82_4_btb_entry = _RAND_43[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_82_4_btb_bht_history = _RAND_44[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {2{`RANDOM}};
  _T_82_4_pc = _RAND_45[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_82_4_data = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_82_4_xcpt_pf_inst = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_82_4_xcpt_ae_inst = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_82_4_replay = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  ShiftQueue_state = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ShiftQueue_cov[initvar] = _RAND_51[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  ShiftQueue_covSum = _RAND_52[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      _T_60_0 <= 1'h0;
    end else if (reset) begin
      _T_60_0 <= 1'h0;
    end else if (io_deq_ready) begin
      _T_60_0 <= _T_94;
    end else begin
      _T_60_0 <= _T_106;
    end
    if (metaReset) begin
      _T_60_1 <= 1'h0;
    end else if (reset) begin
      _T_60_1 <= 1'h0;
    end else if (io_deq_ready) begin
      _T_60_1 <= _T_112;
    end else begin
      _T_60_1 <= _T_124;
    end
    if (metaReset) begin
      _T_60_2 <= 1'h0;
    end else if (reset) begin
      _T_60_2 <= 1'h0;
    end else if (io_deq_ready) begin
      _T_60_2 <= _T_130;
    end else begin
      _T_60_2 <= _T_142;
    end
    if (metaReset) begin
      _T_60_3 <= 1'h0;
    end else if (reset) begin
      _T_60_3 <= 1'h0;
    end else if (io_deq_ready) begin
      _T_60_3 <= _T_148;
    end else begin
      _T_60_3 <= _T_160;
    end
    if (metaReset) begin
      _T_60_4 <= 1'h0;
    end else if (reset) begin
      _T_60_4 <= 1'h0;
    end else if (io_deq_ready) begin
      _T_60_4 <= _T_164;
    end else begin
      _T_60_4 <= _T_177;
    end
    if (metaReset) begin
      _T_82_0_btb_taken <= 1'h0;
    end else if (_T_99) begin
      if (_T_60_1) begin
        _T_82_0_btb_taken <= _T_82_1_btb_taken;
      end else begin
        _T_82_0_btb_taken <= io_enq_bits_btb_taken;
      end
    end
    if (metaReset) begin
      _T_82_0_btb_bridx <= 1'h0;
    end else if (_T_99) begin
      if (_T_60_1) begin
        _T_82_0_btb_bridx <= _T_82_1_btb_bridx;
      end else begin
        _T_82_0_btb_bridx <= io_enq_bits_btb_bridx;
      end
    end
    if (metaReset) begin
      _T_82_0_btb_entry <= 5'h0;
    end else if (_T_99) begin
      if (_T_60_1) begin
        _T_82_0_btb_entry <= _T_82_1_btb_entry;
      end else begin
        _T_82_0_btb_entry <= io_enq_bits_btb_entry;
      end
    end
    if (metaReset) begin
      _T_82_0_btb_bht_history <= 8'h0;
    end else if (_T_99) begin
      if (_T_60_1) begin
        _T_82_0_btb_bht_history <= _T_82_1_btb_bht_history;
      end else begin
        _T_82_0_btb_bht_history <= io_enq_bits_btb_bht_history;
      end
    end
    if (metaReset) begin
      _T_82_0_pc <= 40'h0;
    end else if (_T_99) begin
      if (_T_60_1) begin
        _T_82_0_pc <= _T_82_1_pc;
      end else begin
        _T_82_0_pc <= io_enq_bits_pc;
      end
    end
    if (metaReset) begin
      _T_82_0_data <= 32'h0;
    end else if (_T_99) begin
      if (_T_60_1) begin
        _T_82_0_data <= _T_82_1_data;
      end else begin
        _T_82_0_data <= io_enq_bits_data;
      end
    end
    if (metaReset) begin
      _T_82_0_xcpt_pf_inst <= 1'h0;
    end else if (_T_99) begin
      if (_T_60_1) begin
        _T_82_0_xcpt_pf_inst <= _T_82_1_xcpt_pf_inst;
      end else begin
        _T_82_0_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
      end
    end
    if (metaReset) begin
      _T_82_0_xcpt_ae_inst <= 1'h0;
    end else if (_T_99) begin
      if (_T_60_1) begin
        _T_82_0_xcpt_ae_inst <= _T_82_1_xcpt_ae_inst;
      end else begin
        _T_82_0_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
      end
    end
    if (metaReset) begin
      _T_82_0_replay <= 1'h0;
    end else if (_T_99) begin
      if (_T_60_1) begin
        _T_82_0_replay <= _T_82_1_replay;
      end else begin
        _T_82_0_replay <= io_enq_bits_replay;
      end
    end
    if (metaReset) begin
      _T_82_1_btb_taken <= 1'h0;
    end else if (_T_117) begin
      if (_T_60_2) begin
        _T_82_1_btb_taken <= _T_82_2_btb_taken;
      end else begin
        _T_82_1_btb_taken <= io_enq_bits_btb_taken;
      end
    end
    if (metaReset) begin
      _T_82_1_btb_bridx <= 1'h0;
    end else if (_T_117) begin
      if (_T_60_2) begin
        _T_82_1_btb_bridx <= _T_82_2_btb_bridx;
      end else begin
        _T_82_1_btb_bridx <= io_enq_bits_btb_bridx;
      end
    end
    if (metaReset) begin
      _T_82_1_btb_entry <= 5'h0;
    end else if (_T_117) begin
      if (_T_60_2) begin
        _T_82_1_btb_entry <= _T_82_2_btb_entry;
      end else begin
        _T_82_1_btb_entry <= io_enq_bits_btb_entry;
      end
    end
    if (metaReset) begin
      _T_82_1_btb_bht_history <= 8'h0;
    end else if (_T_117) begin
      if (_T_60_2) begin
        _T_82_1_btb_bht_history <= _T_82_2_btb_bht_history;
      end else begin
        _T_82_1_btb_bht_history <= io_enq_bits_btb_bht_history;
      end
    end
    if (metaReset) begin
      _T_82_1_pc <= 40'h0;
    end else if (_T_117) begin
      if (_T_60_2) begin
        _T_82_1_pc <= _T_82_2_pc;
      end else begin
        _T_82_1_pc <= io_enq_bits_pc;
      end
    end
    if (metaReset) begin
      _T_82_1_data <= 32'h0;
    end else if (_T_117) begin
      if (_T_60_2) begin
        _T_82_1_data <= _T_82_2_data;
      end else begin
        _T_82_1_data <= io_enq_bits_data;
      end
    end
    if (metaReset) begin
      _T_82_1_xcpt_pf_inst <= 1'h0;
    end else if (_T_117) begin
      if (_T_60_2) begin
        _T_82_1_xcpt_pf_inst <= _T_82_2_xcpt_pf_inst;
      end else begin
        _T_82_1_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
      end
    end
    if (metaReset) begin
      _T_82_1_xcpt_ae_inst <= 1'h0;
    end else if (_T_117) begin
      if (_T_60_2) begin
        _T_82_1_xcpt_ae_inst <= _T_82_2_xcpt_ae_inst;
      end else begin
        _T_82_1_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
      end
    end
    if (metaReset) begin
      _T_82_1_replay <= 1'h0;
    end else if (_T_117) begin
      if (_T_60_2) begin
        _T_82_1_replay <= _T_82_2_replay;
      end else begin
        _T_82_1_replay <= io_enq_bits_replay;
      end
    end
    if (metaReset) begin
      _T_82_2_btb_taken <= 1'h0;
    end else if (_T_135) begin
      if (_T_60_3) begin
        _T_82_2_btb_taken <= _T_82_3_btb_taken;
      end else begin
        _T_82_2_btb_taken <= io_enq_bits_btb_taken;
      end
    end
    if (metaReset) begin
      _T_82_2_btb_bridx <= 1'h0;
    end else if (_T_135) begin
      if (_T_60_3) begin
        _T_82_2_btb_bridx <= _T_82_3_btb_bridx;
      end else begin
        _T_82_2_btb_bridx <= io_enq_bits_btb_bridx;
      end
    end
    if (metaReset) begin
      _T_82_2_btb_entry <= 5'h0;
    end else if (_T_135) begin
      if (_T_60_3) begin
        _T_82_2_btb_entry <= _T_82_3_btb_entry;
      end else begin
        _T_82_2_btb_entry <= io_enq_bits_btb_entry;
      end
    end
    if (metaReset) begin
      _T_82_2_btb_bht_history <= 8'h0;
    end else if (_T_135) begin
      if (_T_60_3) begin
        _T_82_2_btb_bht_history <= _T_82_3_btb_bht_history;
      end else begin
        _T_82_2_btb_bht_history <= io_enq_bits_btb_bht_history;
      end
    end
    if (metaReset) begin
      _T_82_2_pc <= 40'h0;
    end else if (_T_135) begin
      if (_T_60_3) begin
        _T_82_2_pc <= _T_82_3_pc;
      end else begin
        _T_82_2_pc <= io_enq_bits_pc;
      end
    end
    if (metaReset) begin
      _T_82_2_data <= 32'h0;
    end else if (_T_135) begin
      if (_T_60_3) begin
        _T_82_2_data <= _T_82_3_data;
      end else begin
        _T_82_2_data <= io_enq_bits_data;
      end
    end
    if (metaReset) begin
      _T_82_2_xcpt_pf_inst <= 1'h0;
    end else if (_T_135) begin
      if (_T_60_3) begin
        _T_82_2_xcpt_pf_inst <= _T_82_3_xcpt_pf_inst;
      end else begin
        _T_82_2_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
      end
    end
    if (metaReset) begin
      _T_82_2_xcpt_ae_inst <= 1'h0;
    end else if (_T_135) begin
      if (_T_60_3) begin
        _T_82_2_xcpt_ae_inst <= _T_82_3_xcpt_ae_inst;
      end else begin
        _T_82_2_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
      end
    end
    if (metaReset) begin
      _T_82_2_replay <= 1'h0;
    end else if (_T_135) begin
      if (_T_60_3) begin
        _T_82_2_replay <= _T_82_3_replay;
      end else begin
        _T_82_2_replay <= io_enq_bits_replay;
      end
    end
    if (metaReset) begin
      _T_82_3_btb_taken <= 1'h0;
    end else if (_T_153) begin
      if (_T_60_4) begin
        _T_82_3_btb_taken <= _T_82_4_btb_taken;
      end else begin
        _T_82_3_btb_taken <= io_enq_bits_btb_taken;
      end
    end
    if (metaReset) begin
      _T_82_3_btb_bridx <= 1'h0;
    end else if (_T_153) begin
      if (_T_60_4) begin
        _T_82_3_btb_bridx <= _T_82_4_btb_bridx;
      end else begin
        _T_82_3_btb_bridx <= io_enq_bits_btb_bridx;
      end
    end
    if (metaReset) begin
      _T_82_3_btb_entry <= 5'h0;
    end else if (_T_153) begin
      if (_T_60_4) begin
        _T_82_3_btb_entry <= _T_82_4_btb_entry;
      end else begin
        _T_82_3_btb_entry <= io_enq_bits_btb_entry;
      end
    end
    if (metaReset) begin
      _T_82_3_btb_bht_history <= 8'h0;
    end else if (_T_153) begin
      if (_T_60_4) begin
        _T_82_3_btb_bht_history <= _T_82_4_btb_bht_history;
      end else begin
        _T_82_3_btb_bht_history <= io_enq_bits_btb_bht_history;
      end
    end
    if (metaReset) begin
      _T_82_3_pc <= 40'h0;
    end else if (_T_153) begin
      if (_T_60_4) begin
        _T_82_3_pc <= _T_82_4_pc;
      end else begin
        _T_82_3_pc <= io_enq_bits_pc;
      end
    end
    if (metaReset) begin
      _T_82_3_data <= 32'h0;
    end else if (_T_153) begin
      if (_T_60_4) begin
        _T_82_3_data <= _T_82_4_data;
      end else begin
        _T_82_3_data <= io_enq_bits_data;
      end
    end
    if (metaReset) begin
      _T_82_3_xcpt_pf_inst <= 1'h0;
    end else if (_T_153) begin
      if (_T_60_4) begin
        _T_82_3_xcpt_pf_inst <= _T_82_4_xcpt_pf_inst;
      end else begin
        _T_82_3_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
      end
    end
    if (metaReset) begin
      _T_82_3_xcpt_ae_inst <= 1'h0;
    end else if (_T_153) begin
      if (_T_60_4) begin
        _T_82_3_xcpt_ae_inst <= _T_82_4_xcpt_ae_inst;
      end else begin
        _T_82_3_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
      end
    end
    if (metaReset) begin
      _T_82_3_replay <= 1'h0;
    end else if (_T_153) begin
      if (_T_60_4) begin
        _T_82_3_replay <= _T_82_4_replay;
      end else begin
        _T_82_3_replay <= io_enq_bits_replay;
      end
    end
    if (metaReset) begin
      _T_82_4_btb_taken <= 1'h0;
    end else if (_T_170) begin
      _T_82_4_btb_taken <= io_enq_bits_btb_taken;
    end
    if (metaReset) begin
      _T_82_4_btb_bridx <= 1'h0;
    end else if (_T_170) begin
      _T_82_4_btb_bridx <= io_enq_bits_btb_bridx;
    end
    if (metaReset) begin
      _T_82_4_btb_entry <= 5'h0;
    end else if (_T_170) begin
      _T_82_4_btb_entry <= io_enq_bits_btb_entry;
    end
    if (metaReset) begin
      _T_82_4_btb_bht_history <= 8'h0;
    end else if (_T_170) begin
      _T_82_4_btb_bht_history <= io_enq_bits_btb_bht_history;
    end
    if (metaReset) begin
      _T_82_4_pc <= 40'h0;
    end else if (_T_170) begin
      _T_82_4_pc <= io_enq_bits_pc;
    end
    if (metaReset) begin
      _T_82_4_data <= 32'h0;
    end else if (_T_170) begin
      _T_82_4_data <= io_enq_bits_data;
    end
    if (metaReset) begin
      _T_82_4_xcpt_pf_inst <= 1'h0;
    end else if (_T_170) begin
      _T_82_4_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
    end
    if (metaReset) begin
      _T_82_4_xcpt_ae_inst <= 1'h0;
    end else if (_T_170) begin
      _T_82_4_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
    end
    if (metaReset) begin
      _T_82_4_replay <= 1'h0;
    end else if (_T_170) begin
      _T_82_4_replay <= io_enq_bits_replay;
    end
    ShiftQueue_state <= ShiftQueue_xor0;
    if (!(ShiftQueue_cov_read_data)) begin
      ShiftQueue_covSum <= ShiftQueue_covSum + 1'h1;
    end
  end
  always @(posedge clock) begin
    if(ShiftQueue_cov_write_en & ShiftQueue_cov_write_mask) begin
      ShiftQueue_cov[ShiftQueue_cov_write_addr] <= ShiftQueue_cov_write_data; // @[Coverage map for ShiftQueue]
    end
  end
endmodule
module TLB_1(
  input         clock,
  input         reset,
  output        io_req_ready,
  input         io_req_valid,
  input  [39:0] io_req_bits_vaddr,
  output        io_resp_miss,
  output [31:0] io_resp_paddr,
  output        io_resp_pf_inst,
  output        io_resp_ae_inst,
  output        io_resp_cacheable,
  input         io_sfence_valid,
  input         io_sfence_bits_rs1,
  input         io_sfence_bits_rs2,
  input  [38:0] io_sfence_bits_addr,
  input         io_ptw_req_ready,
  output        io_ptw_req_valid,
  output        io_ptw_req_bits_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  input         io_ptw_resp_valid,
  input         io_ptw_resp_bits_ae,
  input  [53:0] io_ptw_resp_bits_pte_ppn,
  input         io_ptw_resp_bits_pte_d,
  input         io_ptw_resp_bits_pte_a,
  input         io_ptw_resp_bits_pte_g,
  input         io_ptw_resp_bits_pte_u,
  input         io_ptw_resp_bits_pte_x,
  input         io_ptw_resp_bits_pte_w,
  input         io_ptw_resp_bits_pte_r,
  input         io_ptw_resp_bits_pte_v,
  input  [1:0]  io_ptw_resp_bits_level,
  input         io_ptw_resp_bits_homogeneous,
  input  [3:0]  io_ptw_ptbr_mode,
  input  [1:0]  io_ptw_status_prv,
  input         io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
  input         io_ptw_pmp_0_cfg_w,
  input         io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr,
  input  [31:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
  input         io_ptw_pmp_1_cfg_w,
  input         io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr,
  input  [31:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
  input         io_ptw_pmp_2_cfg_w,
  input         io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr,
  input  [31:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
  input         io_ptw_pmp_3_cfg_w,
  input         io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr,
  input  [31:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
  input         io_ptw_pmp_4_cfg_w,
  input         io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr,
  input  [31:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
  input         io_ptw_pmp_5_cfg_w,
  input         io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr,
  input  [31:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
  input         io_ptw_pmp_6_cfg_w,
  input         io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr,
  input  [31:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
  input         io_ptw_pmp_7_cfg_w,
  input         io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr,
  input  [31:0] io_ptw_pmp_7_mask,
  input  [26:0] io_ptw_vpoffset_bits_value,
  input         io_kill,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [1:0] pmp_io_prv; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_0_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_0_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_0_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_0_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_0_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_0_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_0_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_1_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_1_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_1_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_1_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_1_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_1_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_1_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_2_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_2_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_2_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_2_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_2_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_2_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_2_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_3_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_3_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_3_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_3_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_3_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_3_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_3_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_4_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_4_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_4_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_4_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_4_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_4_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_4_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_5_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_5_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_5_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_5_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_5_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_5_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_5_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_6_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_6_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_6_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_6_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_6_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_6_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_6_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_7_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_7_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_7_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_7_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_7_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_7_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_7_mask; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_addr; // @[TLB.scala 190:19]
  wire  pmp_io_r; // @[TLB.scala 190:19]
  wire  pmp_io_w; // @[TLB.scala 190:19]
  wire  pmp_io_x; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_covSum; // @[TLB.scala 190:19]
  wire  pmp_metaAssert; // @[TLB.scala 190:19]
  reg [26:0] sectored_entries_0_tag; // @[TLB.scala 163:29]
  reg [31:0] _RAND_0;
  reg [33:0] sectored_entries_0_data_0; // @[TLB.scala 163:29]
  reg [63:0] _RAND_1;
  reg [33:0] sectored_entries_0_data_1; // @[TLB.scala 163:29]
  reg [63:0] _RAND_2;
  reg [33:0] sectored_entries_0_data_2; // @[TLB.scala 163:29]
  reg [63:0] _RAND_3;
  reg [33:0] sectored_entries_0_data_3; // @[TLB.scala 163:29]
  reg [63:0] _RAND_4;
  reg  sectored_entries_0_valid_0; // @[TLB.scala 163:29]
  reg [31:0] _RAND_5;
  reg  sectored_entries_0_valid_1; // @[TLB.scala 163:29]
  reg [31:0] _RAND_6;
  reg  sectored_entries_0_valid_2; // @[TLB.scala 163:29]
  reg [31:0] _RAND_7;
  reg  sectored_entries_0_valid_3; // @[TLB.scala 163:29]
  reg [31:0] _RAND_8;
  reg [26:0] sectored_entries_1_tag; // @[TLB.scala 163:29]
  reg [31:0] _RAND_9;
  reg [33:0] sectored_entries_1_data_0; // @[TLB.scala 163:29]
  reg [63:0] _RAND_10;
  reg [33:0] sectored_entries_1_data_1; // @[TLB.scala 163:29]
  reg [63:0] _RAND_11;
  reg [33:0] sectored_entries_1_data_2; // @[TLB.scala 163:29]
  reg [63:0] _RAND_12;
  reg [33:0] sectored_entries_1_data_3; // @[TLB.scala 163:29]
  reg [63:0] _RAND_13;
  reg  sectored_entries_1_valid_0; // @[TLB.scala 163:29]
  reg [31:0] _RAND_14;
  reg  sectored_entries_1_valid_1; // @[TLB.scala 163:29]
  reg [31:0] _RAND_15;
  reg  sectored_entries_1_valid_2; // @[TLB.scala 163:29]
  reg [31:0] _RAND_16;
  reg  sectored_entries_1_valid_3; // @[TLB.scala 163:29]
  reg [31:0] _RAND_17;
  reg [26:0] sectored_entries_2_tag; // @[TLB.scala 163:29]
  reg [31:0] _RAND_18;
  reg [33:0] sectored_entries_2_data_0; // @[TLB.scala 163:29]
  reg [63:0] _RAND_19;
  reg [33:0] sectored_entries_2_data_1; // @[TLB.scala 163:29]
  reg [63:0] _RAND_20;
  reg [33:0] sectored_entries_2_data_2; // @[TLB.scala 163:29]
  reg [63:0] _RAND_21;
  reg [33:0] sectored_entries_2_data_3; // @[TLB.scala 163:29]
  reg [63:0] _RAND_22;
  reg  sectored_entries_2_valid_0; // @[TLB.scala 163:29]
  reg [31:0] _RAND_23;
  reg  sectored_entries_2_valid_1; // @[TLB.scala 163:29]
  reg [31:0] _RAND_24;
  reg  sectored_entries_2_valid_2; // @[TLB.scala 163:29]
  reg [31:0] _RAND_25;
  reg  sectored_entries_2_valid_3; // @[TLB.scala 163:29]
  reg [31:0] _RAND_26;
  reg [26:0] sectored_entries_3_tag; // @[TLB.scala 163:29]
  reg [31:0] _RAND_27;
  reg [33:0] sectored_entries_3_data_0; // @[TLB.scala 163:29]
  reg [63:0] _RAND_28;
  reg [33:0] sectored_entries_3_data_1; // @[TLB.scala 163:29]
  reg [63:0] _RAND_29;
  reg [33:0] sectored_entries_3_data_2; // @[TLB.scala 163:29]
  reg [63:0] _RAND_30;
  reg [33:0] sectored_entries_3_data_3; // @[TLB.scala 163:29]
  reg [63:0] _RAND_31;
  reg  sectored_entries_3_valid_0; // @[TLB.scala 163:29]
  reg [31:0] _RAND_32;
  reg  sectored_entries_3_valid_1; // @[TLB.scala 163:29]
  reg [31:0] _RAND_33;
  reg  sectored_entries_3_valid_2; // @[TLB.scala 163:29]
  reg [31:0] _RAND_34;
  reg  sectored_entries_3_valid_3; // @[TLB.scala 163:29]
  reg [31:0] _RAND_35;
  reg [26:0] sectored_entries_4_tag; // @[TLB.scala 163:29]
  reg [31:0] _RAND_36;
  reg [33:0] sectored_entries_4_data_0; // @[TLB.scala 163:29]
  reg [63:0] _RAND_37;
  reg [33:0] sectored_entries_4_data_1; // @[TLB.scala 163:29]
  reg [63:0] _RAND_38;
  reg [33:0] sectored_entries_4_data_2; // @[TLB.scala 163:29]
  reg [63:0] _RAND_39;
  reg [33:0] sectored_entries_4_data_3; // @[TLB.scala 163:29]
  reg [63:0] _RAND_40;
  reg  sectored_entries_4_valid_0; // @[TLB.scala 163:29]
  reg [31:0] _RAND_41;
  reg  sectored_entries_4_valid_1; // @[TLB.scala 163:29]
  reg [31:0] _RAND_42;
  reg  sectored_entries_4_valid_2; // @[TLB.scala 163:29]
  reg [31:0] _RAND_43;
  reg  sectored_entries_4_valid_3; // @[TLB.scala 163:29]
  reg [31:0] _RAND_44;
  reg [26:0] sectored_entries_5_tag; // @[TLB.scala 163:29]
  reg [31:0] _RAND_45;
  reg [33:0] sectored_entries_5_data_0; // @[TLB.scala 163:29]
  reg [63:0] _RAND_46;
  reg [33:0] sectored_entries_5_data_1; // @[TLB.scala 163:29]
  reg [63:0] _RAND_47;
  reg [33:0] sectored_entries_5_data_2; // @[TLB.scala 163:29]
  reg [63:0] _RAND_48;
  reg [33:0] sectored_entries_5_data_3; // @[TLB.scala 163:29]
  reg [63:0] _RAND_49;
  reg  sectored_entries_5_valid_0; // @[TLB.scala 163:29]
  reg [31:0] _RAND_50;
  reg  sectored_entries_5_valid_1; // @[TLB.scala 163:29]
  reg [31:0] _RAND_51;
  reg  sectored_entries_5_valid_2; // @[TLB.scala 163:29]
  reg [31:0] _RAND_52;
  reg  sectored_entries_5_valid_3; // @[TLB.scala 163:29]
  reg [31:0] _RAND_53;
  reg [26:0] sectored_entries_6_tag; // @[TLB.scala 163:29]
  reg [31:0] _RAND_54;
  reg [33:0] sectored_entries_6_data_0; // @[TLB.scala 163:29]
  reg [63:0] _RAND_55;
  reg [33:0] sectored_entries_6_data_1; // @[TLB.scala 163:29]
  reg [63:0] _RAND_56;
  reg [33:0] sectored_entries_6_data_2; // @[TLB.scala 163:29]
  reg [63:0] _RAND_57;
  reg [33:0] sectored_entries_6_data_3; // @[TLB.scala 163:29]
  reg [63:0] _RAND_58;
  reg  sectored_entries_6_valid_0; // @[TLB.scala 163:29]
  reg [31:0] _RAND_59;
  reg  sectored_entries_6_valid_1; // @[TLB.scala 163:29]
  reg [31:0] _RAND_60;
  reg  sectored_entries_6_valid_2; // @[TLB.scala 163:29]
  reg [31:0] _RAND_61;
  reg  sectored_entries_6_valid_3; // @[TLB.scala 163:29]
  reg [31:0] _RAND_62;
  reg [26:0] sectored_entries_7_tag; // @[TLB.scala 163:29]
  reg [31:0] _RAND_63;
  reg [33:0] sectored_entries_7_data_0; // @[TLB.scala 163:29]
  reg [63:0] _RAND_64;
  reg [33:0] sectored_entries_7_data_1; // @[TLB.scala 163:29]
  reg [63:0] _RAND_65;
  reg [33:0] sectored_entries_7_data_2; // @[TLB.scala 163:29]
  reg [63:0] _RAND_66;
  reg [33:0] sectored_entries_7_data_3; // @[TLB.scala 163:29]
  reg [63:0] _RAND_67;
  reg  sectored_entries_7_valid_0; // @[TLB.scala 163:29]
  reg [31:0] _RAND_68;
  reg  sectored_entries_7_valid_1; // @[TLB.scala 163:29]
  reg [31:0] _RAND_69;
  reg  sectored_entries_7_valid_2; // @[TLB.scala 163:29]
  reg [31:0] _RAND_70;
  reg  sectored_entries_7_valid_3; // @[TLB.scala 163:29]
  reg [31:0] _RAND_71;
  reg [1:0] superpage_entries_0_level; // @[TLB.scala 164:30]
  reg [31:0] _RAND_72;
  reg [26:0] superpage_entries_0_tag; // @[TLB.scala 164:30]
  reg [31:0] _RAND_73;
  reg [33:0] superpage_entries_0_data_0; // @[TLB.scala 164:30]
  reg [63:0] _RAND_74;
  reg  superpage_entries_0_valid_0; // @[TLB.scala 164:30]
  reg [31:0] _RAND_75;
  reg [1:0] superpage_entries_1_level; // @[TLB.scala 164:30]
  reg [31:0] _RAND_76;
  reg [26:0] superpage_entries_1_tag; // @[TLB.scala 164:30]
  reg [31:0] _RAND_77;
  reg [33:0] superpage_entries_1_data_0; // @[TLB.scala 164:30]
  reg [63:0] _RAND_78;
  reg  superpage_entries_1_valid_0; // @[TLB.scala 164:30]
  reg [31:0] _RAND_79;
  reg [1:0] superpage_entries_2_level; // @[TLB.scala 164:30]
  reg [31:0] _RAND_80;
  reg [26:0] superpage_entries_2_tag; // @[TLB.scala 164:30]
  reg [31:0] _RAND_81;
  reg [33:0] superpage_entries_2_data_0; // @[TLB.scala 164:30]
  reg [63:0] _RAND_82;
  reg  superpage_entries_2_valid_0; // @[TLB.scala 164:30]
  reg [31:0] _RAND_83;
  reg [1:0] superpage_entries_3_level; // @[TLB.scala 164:30]
  reg [31:0] _RAND_84;
  reg [26:0] superpage_entries_3_tag; // @[TLB.scala 164:30]
  reg [31:0] _RAND_85;
  reg [33:0] superpage_entries_3_data_0; // @[TLB.scala 164:30]
  reg [63:0] _RAND_86;
  reg  superpage_entries_3_valid_0; // @[TLB.scala 164:30]
  reg [31:0] _RAND_87;
  reg [1:0] special_entry_level; // @[TLB.scala 165:56]
  reg [31:0] _RAND_88;
  reg [26:0] special_entry_tag; // @[TLB.scala 165:56]
  reg [31:0] _RAND_89;
  reg [33:0] special_entry_data_0; // @[TLB.scala 165:56]
  reg [63:0] _RAND_90;
  reg  special_entry_valid_0; // @[TLB.scala 165:56]
  reg [31:0] _RAND_91;
  reg [1:0] state; // @[TLB.scala 170:18]
  reg [31:0] _RAND_92;
  reg [26:0] r_refill_tag; // @[TLB.scala 171:25]
  reg [31:0] _RAND_93;
  reg [1:0] r_superpage_repl_addr; // @[TLB.scala 172:34]
  reg [31:0] _RAND_94;
  reg [2:0] r_sectored_repl_addr; // @[TLB.scala 173:33]
  reg [31:0] _RAND_95;
  reg [2:0] r_sectored_hit_addr; // @[TLB.scala 174:32]
  reg [31:0] _RAND_96;
  reg  r_sectored_hit; // @[TLB.scala 175:27]
  reg [31:0] _RAND_97;
  wire  priv_s; // @[TLB.scala 178:20]
  wire  priv_uses_vm; // @[TLB.scala 179:27]
  wire  vm_enabled; // @[TLB.scala 180:83]
  wire [26:0] vpn; // @[TLB.scala 183:30]
  wire [19:0] refill_ppn; // @[TLB.scala 184:44]
  wire  _T_324; // @[package.scala 14:47]
  wire  _T_325; // @[package.scala 14:47]
  wire  invalidate_refill; // @[package.scala 14:62]
  wire  _T_348; // @[TLB.scala 123:30]
  wire [26:0] _T_350; // @[TLB.scala 124:30]
  wire [26:0] _GEN_954; // @[TLB.scala 124:49]
  wire [26:0] _T_351; // @[TLB.scala 124:49]
  wire  _T_354; // @[TLB.scala 123:30]
  wire [26:0] _T_356; // @[TLB.scala 124:30]
  wire [26:0] _T_357; // @[TLB.scala 124:49]
  wire [19:0] _T_359; // @[Cat.scala 30:58]
  wire [27:0] _T_361; // @[TLB.scala 188:20]
  wire [27:0] mpu_ppn; // @[TLB.scala 187:20]
  wire [39:0] mpu_physaddr; // @[Cat.scala 30:58]
  wire [39:0] _T_366; // @[Parameters.scala 121:31]
  wire [40:0] _T_367; // @[Parameters.scala 121:49]
  wire [40:0] _T_369; // @[Parameters.scala 121:52]
  wire  _T_370; // @[Parameters.scala 121:67]
  wire [39:0] _T_371; // @[Parameters.scala 121:31]
  wire [40:0] _T_372; // @[Parameters.scala 121:49]
  wire [40:0] _T_374; // @[Parameters.scala 121:52]
  wire  _T_375; // @[Parameters.scala 121:67]
  wire [39:0] _T_376; // @[Parameters.scala 121:31]
  wire [40:0] _T_377; // @[Parameters.scala 121:49]
  wire [40:0] _T_379; // @[Parameters.scala 121:52]
  wire  _T_380; // @[Parameters.scala 121:67]
  wire [40:0] _T_382; // @[Parameters.scala 121:49]
  wire [40:0] _T_384; // @[Parameters.scala 121:52]
  wire  _T_385; // @[Parameters.scala 121:67]
  wire [39:0] _T_386; // @[Parameters.scala 121:31]
  wire [40:0] _T_387; // @[Parameters.scala 121:49]
  wire [40:0] _T_389; // @[Parameters.scala 121:52]
  wire  _T_390; // @[Parameters.scala 121:67]
  wire [39:0] _T_391; // @[Parameters.scala 121:31]
  wire [40:0] _T_392; // @[Parameters.scala 121:49]
  wire [40:0] _T_394; // @[Parameters.scala 121:52]
  wire  _T_395; // @[Parameters.scala 121:67]
  wire [39:0] _T_396; // @[Parameters.scala 121:31]
  wire [40:0] _T_397; // @[Parameters.scala 121:49]
  wire [40:0] _T_399; // @[Parameters.scala 121:52]
  wire  _T_400; // @[Parameters.scala 121:67]
  wire  _T_414; // @[TLB.scala 195:67]
  wire  _T_415; // @[TLB.scala 195:67]
  wire  _T_416; // @[TLB.scala 195:67]
  wire  _T_417; // @[TLB.scala 195:67]
  wire  _T_418; // @[TLB.scala 195:67]
  wire  legal_address; // @[TLB.scala 195:67]
  wire [40:0] _T_427; // @[Parameters.scala 121:52]
  wire  _T_428; // @[Parameters.scala 121:67]
  wire  cacheable; // @[TLB.scala 197:19]
  wire [39:0] _T_485; // @[Parameters.scala 121:31]
  wire [40:0] _T_486; // @[Parameters.scala 121:49]
  wire [40:0] _T_488; // @[Parameters.scala 121:52]
  wire  _T_489; // @[Parameters.scala 121:67]
  wire [40:0] _T_507; // @[Parameters.scala 121:52]
  wire  _T_508; // @[Parameters.scala 121:67]
  wire  _T_515; // @[TLBPermissions.scala 81:66]
  wire  prot_r; // @[TLB.scala 200:41]
  wire [40:0] _T_552; // @[Parameters.scala 121:52]
  wire  _T_553; // @[Parameters.scala 121:67]
  wire [39:0] _T_554; // @[Parameters.scala 121:31]
  wire [40:0] _T_555; // @[Parameters.scala 121:49]
  wire [40:0] _T_557; // @[Parameters.scala 121:52]
  wire  _T_558; // @[Parameters.scala 121:67]
  wire  _T_560; // @[Parameters.scala 148:89]
  wire  _T_561; // @[Parameters.scala 148:89]
  wire  _T_568; // @[TLB.scala 197:19]
  wire  prot_w; // @[TLB.scala 201:45]
  wire  _T_603; // @[TLB.scala 197:19]
  wire  prot_al; // @[TLB.scala 202:46]
  wire [40:0] _T_655; // @[Parameters.scala 121:52]
  wire  _T_656; // @[Parameters.scala 121:67]
  wire  _T_667; // @[Parameters.scala 148:89]
  wire  _T_668; // @[Parameters.scala 148:89]
  wire  _T_675; // @[TLB.scala 197:19]
  wire  prot_x; // @[TLB.scala 204:40]
  wire [40:0] _T_701; // @[Parameters.scala 121:52]
  wire  _T_702; // @[Parameters.scala 121:67]
  wire [40:0] _T_706; // @[Parameters.scala 121:52]
  wire  _T_707; // @[Parameters.scala 121:67]
  wire  _T_713; // @[Parameters.scala 148:89]
  wire  _T_714; // @[Parameters.scala 148:89]
  wire  _T_715; // @[Parameters.scala 148:89]
  wire  prot_eff; // @[TLB.scala 197:19]
  wire  _T_722; // @[package.scala 63:59]
  wire  _T_723; // @[package.scala 63:59]
  wire  _T_724; // @[package.scala 63:59]
  wire [26:0] _T_725; // @[TLB.scala 103:43]
  wire  _T_727; // @[TLB.scala 103:68]
  wire  sector_hits_0; // @[TLB.scala 102:42]
  wire  _T_728; // @[package.scala 63:59]
  wire  _T_729; // @[package.scala 63:59]
  wire  _T_730; // @[package.scala 63:59]
  wire [26:0] _T_731; // @[TLB.scala 103:43]
  wire  _T_733; // @[TLB.scala 103:68]
  wire  sector_hits_1; // @[TLB.scala 102:42]
  wire  _T_734; // @[package.scala 63:59]
  wire  _T_735; // @[package.scala 63:59]
  wire  _T_736; // @[package.scala 63:59]
  wire [26:0] _T_737; // @[TLB.scala 103:43]
  wire  _T_739; // @[TLB.scala 103:68]
  wire  sector_hits_2; // @[TLB.scala 102:42]
  wire  _T_740; // @[package.scala 63:59]
  wire  _T_741; // @[package.scala 63:59]
  wire  _T_742; // @[package.scala 63:59]
  wire [26:0] _T_743; // @[TLB.scala 103:43]
  wire  _T_745; // @[TLB.scala 103:68]
  wire  sector_hits_3; // @[TLB.scala 102:42]
  wire  _T_746; // @[package.scala 63:59]
  wire  _T_747; // @[package.scala 63:59]
  wire  _T_748; // @[package.scala 63:59]
  wire [26:0] _T_749; // @[TLB.scala 103:43]
  wire  _T_751; // @[TLB.scala 103:68]
  wire  sector_hits_4; // @[TLB.scala 102:42]
  wire  _T_752; // @[package.scala 63:59]
  wire  _T_753; // @[package.scala 63:59]
  wire  _T_754; // @[package.scala 63:59]
  wire [26:0] _T_755; // @[TLB.scala 103:43]
  wire  _T_757; // @[TLB.scala 103:68]
  wire  sector_hits_5; // @[TLB.scala 102:42]
  wire  _T_758; // @[package.scala 63:59]
  wire  _T_759; // @[package.scala 63:59]
  wire  _T_760; // @[package.scala 63:59]
  wire [26:0] _T_761; // @[TLB.scala 103:43]
  wire  _T_763; // @[TLB.scala 103:68]
  wire  sector_hits_6; // @[TLB.scala 102:42]
  wire  _T_764; // @[package.scala 63:59]
  wire  _T_765; // @[package.scala 63:59]
  wire  _T_766; // @[package.scala 63:59]
  wire [26:0] _T_767; // @[TLB.scala 103:43]
  wire  _T_769; // @[TLB.scala 103:68]
  wire  sector_hits_7; // @[TLB.scala 102:42]
  wire  _T_774; // @[TLB.scala 110:79]
  wire  _T_776; // @[TLB.scala 110:31]
  wire  _T_777; // @[TLB.scala 109:30]
  wire  _T_781; // @[TLB.scala 110:79]
  wire  _T_782; // @[TLB.scala 110:42]
  wire  superpage_hits_0; // @[TLB.scala 110:31]
  wire  _T_794; // @[TLB.scala 110:79]
  wire  _T_796; // @[TLB.scala 110:31]
  wire  _T_797; // @[TLB.scala 109:30]
  wire  _T_801; // @[TLB.scala 110:79]
  wire  _T_802; // @[TLB.scala 110:42]
  wire  superpage_hits_1; // @[TLB.scala 110:31]
  wire  _T_814; // @[TLB.scala 110:79]
  wire  _T_816; // @[TLB.scala 110:31]
  wire  _T_817; // @[TLB.scala 109:30]
  wire  _T_821; // @[TLB.scala 110:79]
  wire  _T_822; // @[TLB.scala 110:42]
  wire  superpage_hits_2; // @[TLB.scala 110:31]
  wire  _T_834; // @[TLB.scala 110:79]
  wire  _T_836; // @[TLB.scala 110:31]
  wire  _T_837; // @[TLB.scala 109:30]
  wire  _T_841; // @[TLB.scala 110:79]
  wire  _T_842; // @[TLB.scala 110:42]
  wire  superpage_hits_3; // @[TLB.scala 110:31]
  wire  _GEN_1; // @[TLB.scala 115:20]
  wire  _GEN_2; // @[TLB.scala 115:20]
  wire  _GEN_3; // @[TLB.scala 115:20]
  wire  _T_854; // @[TLB.scala 115:20]
  wire  hitsVec_0; // @[TLB.scala 209:44]
  wire  _GEN_5; // @[TLB.scala 115:20]
  wire  _GEN_6; // @[TLB.scala 115:20]
  wire  _GEN_7; // @[TLB.scala 115:20]
  wire  _T_859; // @[TLB.scala 115:20]
  wire  hitsVec_1; // @[TLB.scala 209:44]
  wire  _GEN_9; // @[TLB.scala 115:20]
  wire  _GEN_10; // @[TLB.scala 115:20]
  wire  _GEN_11; // @[TLB.scala 115:20]
  wire  _T_864; // @[TLB.scala 115:20]
  wire  hitsVec_2; // @[TLB.scala 209:44]
  wire  _GEN_13; // @[TLB.scala 115:20]
  wire  _GEN_14; // @[TLB.scala 115:20]
  wire  _GEN_15; // @[TLB.scala 115:20]
  wire  _T_869; // @[TLB.scala 115:20]
  wire  hitsVec_3; // @[TLB.scala 209:44]
  wire  _GEN_17; // @[TLB.scala 115:20]
  wire  _GEN_18; // @[TLB.scala 115:20]
  wire  _GEN_19; // @[TLB.scala 115:20]
  wire  _T_874; // @[TLB.scala 115:20]
  wire  hitsVec_4; // @[TLB.scala 209:44]
  wire  _GEN_21; // @[TLB.scala 115:20]
  wire  _GEN_22; // @[TLB.scala 115:20]
  wire  _GEN_23; // @[TLB.scala 115:20]
  wire  _T_879; // @[TLB.scala 115:20]
  wire  hitsVec_5; // @[TLB.scala 209:44]
  wire  _GEN_25; // @[TLB.scala 115:20]
  wire  _GEN_26; // @[TLB.scala 115:20]
  wire  _GEN_27; // @[TLB.scala 115:20]
  wire  _T_884; // @[TLB.scala 115:20]
  wire  hitsVec_6; // @[TLB.scala 209:44]
  wire  _GEN_29; // @[TLB.scala 115:20]
  wire  _GEN_30; // @[TLB.scala 115:20]
  wire  _GEN_31; // @[TLB.scala 115:20]
  wire  _T_889; // @[TLB.scala 115:20]
  wire  hitsVec_7; // @[TLB.scala 209:44]
  wire  hitsVec_8; // @[TLB.scala 209:44]
  wire  hitsVec_9; // @[TLB.scala 209:44]
  wire  hitsVec_10; // @[TLB.scala 209:44]
  wire  hitsVec_11; // @[TLB.scala 209:44]
  wire  _T_978; // @[TLB.scala 110:79]
  wire  _T_980; // @[TLB.scala 110:31]
  wire  _T_985; // @[TLB.scala 110:79]
  wire  _T_986; // @[TLB.scala 110:42]
  wire  _T_987; // @[TLB.scala 110:31]
  wire  _T_992; // @[TLB.scala 110:79]
  wire  _T_993; // @[TLB.scala 110:42]
  wire  _T_994; // @[TLB.scala 110:31]
  wire  hitsVec_12; // @[TLB.scala 209:44]
  wire [5:0] _T_999; // @[Cat.scala 30:58]
  wire [12:0] real_hits; // @[Cat.scala 30:58]
  wire [13:0] hits; // @[Cat.scala 30:58]
  wire [33:0] _GEN_33;
  wire [33:0] _GEN_34;
  wire [33:0] _GEN_35;
  wire [33:0] _GEN_37;
  wire [33:0] _GEN_38;
  wire [33:0] _GEN_39;
  wire [33:0] _GEN_41;
  wire [33:0] _GEN_42;
  wire [33:0] _GEN_43;
  wire [33:0] _GEN_45;
  wire [33:0] _GEN_46;
  wire [33:0] _GEN_47;
  wire [33:0] _GEN_49;
  wire [33:0] _GEN_50;
  wire [33:0] _GEN_51;
  wire [33:0] _GEN_53;
  wire [33:0] _GEN_54;
  wire [33:0] _GEN_55;
  wire [33:0] _GEN_57;
  wire [33:0] _GEN_58;
  wire [33:0] _GEN_59;
  wire [33:0] _GEN_61;
  wire [33:0] _GEN_62;
  wire [33:0] _GEN_63;
  wire [26:0] _T_1199; // @[TLB.scala 124:30]
  wire [26:0] _GEN_956; // @[TLB.scala 124:49]
  wire [26:0] _T_1200; // @[TLB.scala 124:49]
  wire [26:0] _T_1206; // @[TLB.scala 124:49]
  wire [19:0] _T_1208; // @[Cat.scala 30:58]
  wire [26:0] _T_1232; // @[TLB.scala 124:30]
  wire [26:0] _GEN_958; // @[TLB.scala 124:49]
  wire [26:0] _T_1233; // @[TLB.scala 124:49]
  wire [26:0] _T_1239; // @[TLB.scala 124:49]
  wire [19:0] _T_1241; // @[Cat.scala 30:58]
  wire [26:0] _T_1265; // @[TLB.scala 124:30]
  wire [26:0] _GEN_960; // @[TLB.scala 124:49]
  wire [26:0] _T_1266; // @[TLB.scala 124:49]
  wire [26:0] _T_1272; // @[TLB.scala 124:49]
  wire [19:0] _T_1274; // @[Cat.scala 30:58]
  wire [26:0] _T_1298; // @[TLB.scala 124:30]
  wire [26:0] _GEN_962; // @[TLB.scala 124:49]
  wire [26:0] _T_1299; // @[TLB.scala 124:49]
  wire [26:0] _T_1305; // @[TLB.scala 124:49]
  wire [19:0] _T_1307; // @[Cat.scala 30:58]
  wire [19:0] _T_1343; // @[Mux.scala 19:72]
  wire [19:0] _T_1344; // @[Mux.scala 19:72]
  wire [19:0] _T_1345; // @[Mux.scala 19:72]
  wire [19:0] _T_1346; // @[Mux.scala 19:72]
  wire [19:0] _T_1347; // @[Mux.scala 19:72]
  wire [19:0] _T_1348; // @[Mux.scala 19:72]
  wire [19:0] _T_1349; // @[Mux.scala 19:72]
  wire [19:0] _T_1350; // @[Mux.scala 19:72]
  wire [19:0] _T_1351; // @[Mux.scala 19:72]
  wire [19:0] _T_1352; // @[Mux.scala 19:72]
  wire [19:0] _T_1353; // @[Mux.scala 19:72]
  wire [19:0] _T_1354; // @[Mux.scala 19:72]
  wire [19:0] _T_1355; // @[Mux.scala 19:72]
  wire [19:0] _T_1356; // @[Mux.scala 19:72]
  wire [19:0] _T_1357; // @[Mux.scala 19:72]
  wire [19:0] _T_1358; // @[Mux.scala 19:72]
  wire [19:0] _T_1359; // @[Mux.scala 19:72]
  wire [19:0] _T_1360; // @[Mux.scala 19:72]
  wire [19:0] _T_1361; // @[Mux.scala 19:72]
  wire [19:0] _T_1362; // @[Mux.scala 19:72]
  wire [19:0] _T_1363; // @[Mux.scala 19:72]
  wire [19:0] _T_1364; // @[Mux.scala 19:72]
  wire [19:0] _T_1365; // @[Mux.scala 19:72]
  wire [19:0] _T_1366; // @[Mux.scala 19:72]
  wire [19:0] _T_1367; // @[Mux.scala 19:72]
  wire [19:0] _T_1368; // @[Mux.scala 19:72]
  wire [19:0] ppn; // @[Mux.scala 19:72]
  reg [26:0] vpoffset_cfg_value; // @[TLB.scala 215:29]
  reg [31:0] _RAND_98;
  reg [26:0] requestedVPN; // @[TLB.scala 216:25]
  reg [31:0] _RAND_99;
  wire  _T_1385; // @[TLB.scala 224:17]
  wire [53:0] _GEN_966; // @[TLB.scala 227:31]
  wire [53:0] _T_1387; // @[TLB.scala 227:31]
  wire  _T_1391; // @[PTW.scala 77:44]
  wire  _T_1392; // @[PTW.scala 77:38]
  wire  _T_1393; // @[PTW.scala 77:32]
  wire  _T_1394; // @[PTW.scala 77:52]
  wire  _T_1395; // @[PTW.scala 81:35]
  wire  _T_1401; // @[PTW.scala 82:35]
  wire  _T_1402; // @[PTW.scala 82:40]
  wire  _T_1403; // @[TLB.scala 231:55]
  wire  _T_1404; // @[TLB.scala 231:32]
  wire  _T_1405; // @[TLB.scala 231:90]
  wire  _T_1406; // @[TLB.scala 231:64]
  wire  _T_1412; // @[PTW.scala 83:35]
  wire [53:0] _GEN_967; // @[TLB.scala 231:133]
  wire  _T_1413; // @[TLB.scala 231:133]
  wire  _T_1420; // @[TLB.scala 231:120]
  wire  _T_1421; // @[TLB.scala 231:25]
  wire [6:0] _T_1430; // @[TLB.scala 138:26]
  wire [33:0] _T_1438; // @[TLB.scala 138:26]
  wire  _T_1439; // @[TLB.scala 253:40]
  wire  _T_1440; // @[TLB.scala 254:82]
  wire  _GEN_67; // @[TLB.scala 254:89]
  wire  _T_1456; // @[TLB.scala 254:82]
  wire  _GEN_71; // @[TLB.scala 254:89]
  wire  _T_1472; // @[TLB.scala 254:82]
  wire  _GEN_75; // @[TLB.scala 254:89]
  wire  _T_1488; // @[TLB.scala 254:82]
  wire  _GEN_79; // @[TLB.scala 254:89]
  wire [2:0] _T_1504; // @[TLB.scala 258:22]
  wire  _T_1505; // @[TLB.scala 259:65]
  wire  _GEN_81; // @[TLB.scala 260:32]
  wire  _GEN_82; // @[TLB.scala 260:32]
  wire  _GEN_83; // @[TLB.scala 260:32]
  wire  _GEN_84; // @[TLB.scala 260:32]
  wire  _GEN_968; // @[TLB.scala 137:18]
  wire  _GEN_85; // @[TLB.scala 137:18]
  wire  _GEN_969; // @[TLB.scala 137:18]
  wire  _GEN_86; // @[TLB.scala 137:18]
  wire  _GEN_970; // @[TLB.scala 137:18]
  wire  _GEN_87; // @[TLB.scala 137:18]
  wire  _GEN_971; // @[TLB.scala 137:18]
  wire  _GEN_88; // @[TLB.scala 137:18]
  wire  _GEN_93; // @[TLB.scala 259:72]
  wire  _GEN_94; // @[TLB.scala 259:72]
  wire  _GEN_95; // @[TLB.scala 259:72]
  wire  _GEN_96; // @[TLB.scala 259:72]
  wire  _T_1522; // @[TLB.scala 259:65]
  wire  _GEN_103; // @[TLB.scala 260:32]
  wire  _GEN_104; // @[TLB.scala 260:32]
  wire  _GEN_105; // @[TLB.scala 260:32]
  wire  _GEN_106; // @[TLB.scala 260:32]
  wire  _GEN_107; // @[TLB.scala 137:18]
  wire  _GEN_108; // @[TLB.scala 137:18]
  wire  _GEN_109; // @[TLB.scala 137:18]
  wire  _GEN_110; // @[TLB.scala 137:18]
  wire  _GEN_115; // @[TLB.scala 259:72]
  wire  _GEN_116; // @[TLB.scala 259:72]
  wire  _GEN_117; // @[TLB.scala 259:72]
  wire  _GEN_118; // @[TLB.scala 259:72]
  wire  _T_1539; // @[TLB.scala 259:65]
  wire  _GEN_125; // @[TLB.scala 260:32]
  wire  _GEN_126; // @[TLB.scala 260:32]
  wire  _GEN_127; // @[TLB.scala 260:32]
  wire  _GEN_128; // @[TLB.scala 260:32]
  wire  _GEN_129; // @[TLB.scala 137:18]
  wire  _GEN_130; // @[TLB.scala 137:18]
  wire  _GEN_131; // @[TLB.scala 137:18]
  wire  _GEN_132; // @[TLB.scala 137:18]
  wire  _GEN_137; // @[TLB.scala 259:72]
  wire  _GEN_138; // @[TLB.scala 259:72]
  wire  _GEN_139; // @[TLB.scala 259:72]
  wire  _GEN_140; // @[TLB.scala 259:72]
  wire  _T_1556; // @[TLB.scala 259:65]
  wire  _GEN_147; // @[TLB.scala 260:32]
  wire  _GEN_148; // @[TLB.scala 260:32]
  wire  _GEN_149; // @[TLB.scala 260:32]
  wire  _GEN_150; // @[TLB.scala 260:32]
  wire  _GEN_151; // @[TLB.scala 137:18]
  wire  _GEN_152; // @[TLB.scala 137:18]
  wire  _GEN_153; // @[TLB.scala 137:18]
  wire  _GEN_154; // @[TLB.scala 137:18]
  wire  _GEN_159; // @[TLB.scala 259:72]
  wire  _GEN_160; // @[TLB.scala 259:72]
  wire  _GEN_161; // @[TLB.scala 259:72]
  wire  _GEN_162; // @[TLB.scala 259:72]
  wire  _T_1573; // @[TLB.scala 259:65]
  wire  _GEN_169; // @[TLB.scala 260:32]
  wire  _GEN_170; // @[TLB.scala 260:32]
  wire  _GEN_171; // @[TLB.scala 260:32]
  wire  _GEN_172; // @[TLB.scala 260:32]
  wire  _GEN_173; // @[TLB.scala 137:18]
  wire  _GEN_174; // @[TLB.scala 137:18]
  wire  _GEN_175; // @[TLB.scala 137:18]
  wire  _GEN_176; // @[TLB.scala 137:18]
  wire  _GEN_181; // @[TLB.scala 259:72]
  wire  _GEN_182; // @[TLB.scala 259:72]
  wire  _GEN_183; // @[TLB.scala 259:72]
  wire  _GEN_184; // @[TLB.scala 259:72]
  wire  _T_1590; // @[TLB.scala 259:65]
  wire  _GEN_191; // @[TLB.scala 260:32]
  wire  _GEN_192; // @[TLB.scala 260:32]
  wire  _GEN_193; // @[TLB.scala 260:32]
  wire  _GEN_194; // @[TLB.scala 260:32]
  wire  _GEN_195; // @[TLB.scala 137:18]
  wire  _GEN_196; // @[TLB.scala 137:18]
  wire  _GEN_197; // @[TLB.scala 137:18]
  wire  _GEN_198; // @[TLB.scala 137:18]
  wire  _GEN_203; // @[TLB.scala 259:72]
  wire  _GEN_204; // @[TLB.scala 259:72]
  wire  _GEN_205; // @[TLB.scala 259:72]
  wire  _GEN_206; // @[TLB.scala 259:72]
  wire  _T_1607; // @[TLB.scala 259:65]
  wire  _GEN_213; // @[TLB.scala 260:32]
  wire  _GEN_214; // @[TLB.scala 260:32]
  wire  _GEN_215; // @[TLB.scala 260:32]
  wire  _GEN_216; // @[TLB.scala 260:32]
  wire  _GEN_217; // @[TLB.scala 137:18]
  wire  _GEN_218; // @[TLB.scala 137:18]
  wire  _GEN_219; // @[TLB.scala 137:18]
  wire  _GEN_220; // @[TLB.scala 137:18]
  wire  _GEN_225; // @[TLB.scala 259:72]
  wire  _GEN_226; // @[TLB.scala 259:72]
  wire  _GEN_227; // @[TLB.scala 259:72]
  wire  _GEN_228; // @[TLB.scala 259:72]
  wire  _T_1624; // @[TLB.scala 259:65]
  wire  _GEN_235; // @[TLB.scala 260:32]
  wire  _GEN_236; // @[TLB.scala 260:32]
  wire  _GEN_237; // @[TLB.scala 260:32]
  wire  _GEN_238; // @[TLB.scala 260:32]
  wire  _GEN_239; // @[TLB.scala 137:18]
  wire  _GEN_240; // @[TLB.scala 137:18]
  wire  _GEN_241; // @[TLB.scala 137:18]
  wire  _GEN_242; // @[TLB.scala 137:18]
  wire  _GEN_247; // @[TLB.scala 259:72]
  wire  _GEN_248; // @[TLB.scala 259:72]
  wire  _GEN_249; // @[TLB.scala 259:72]
  wire  _GEN_250; // @[TLB.scala 259:72]
  wire  _GEN_259; // @[TLB.scala 253:54]
  wire  _GEN_263; // @[TLB.scala 253:54]
  wire  _GEN_267; // @[TLB.scala 253:54]
  wire  _GEN_271; // @[TLB.scala 253:54]
  wire  _GEN_273; // @[TLB.scala 253:54]
  wire  _GEN_274; // @[TLB.scala 253:54]
  wire  _GEN_275; // @[TLB.scala 253:54]
  wire  _GEN_276; // @[TLB.scala 253:54]
  wire  _GEN_283; // @[TLB.scala 253:54]
  wire  _GEN_284; // @[TLB.scala 253:54]
  wire  _GEN_285; // @[TLB.scala 253:54]
  wire  _GEN_286; // @[TLB.scala 253:54]
  wire  _GEN_293; // @[TLB.scala 253:54]
  wire  _GEN_294; // @[TLB.scala 253:54]
  wire  _GEN_295; // @[TLB.scala 253:54]
  wire  _GEN_296; // @[TLB.scala 253:54]
  wire  _GEN_303; // @[TLB.scala 253:54]
  wire  _GEN_304; // @[TLB.scala 253:54]
  wire  _GEN_305; // @[TLB.scala 253:54]
  wire  _GEN_306; // @[TLB.scala 253:54]
  wire  _GEN_313; // @[TLB.scala 253:54]
  wire  _GEN_314; // @[TLB.scala 253:54]
  wire  _GEN_315; // @[TLB.scala 253:54]
  wire  _GEN_316; // @[TLB.scala 253:54]
  wire  _GEN_323; // @[TLB.scala 253:54]
  wire  _GEN_324; // @[TLB.scala 253:54]
  wire  _GEN_325; // @[TLB.scala 253:54]
  wire  _GEN_326; // @[TLB.scala 253:54]
  wire  _GEN_333; // @[TLB.scala 253:54]
  wire  _GEN_334; // @[TLB.scala 253:54]
  wire  _GEN_335; // @[TLB.scala 253:54]
  wire  _GEN_336; // @[TLB.scala 253:54]
  wire  _GEN_343; // @[TLB.scala 253:54]
  wire  _GEN_344; // @[TLB.scala 253:54]
  wire  _GEN_345; // @[TLB.scala 253:54]
  wire  _GEN_346; // @[TLB.scala 253:54]
  wire  _GEN_355; // @[TLB.scala 251:68]
  wire  _GEN_359; // @[TLB.scala 251:68]
  wire  _GEN_363; // @[TLB.scala 251:68]
  wire  _GEN_367; // @[TLB.scala 251:68]
  wire  _GEN_371; // @[TLB.scala 251:68]
  wire  _GEN_373; // @[TLB.scala 251:68]
  wire  _GEN_374; // @[TLB.scala 251:68]
  wire  _GEN_375; // @[TLB.scala 251:68]
  wire  _GEN_376; // @[TLB.scala 251:68]
  wire  _GEN_383; // @[TLB.scala 251:68]
  wire  _GEN_384; // @[TLB.scala 251:68]
  wire  _GEN_385; // @[TLB.scala 251:68]
  wire  _GEN_386; // @[TLB.scala 251:68]
  wire  _GEN_393; // @[TLB.scala 251:68]
  wire  _GEN_394; // @[TLB.scala 251:68]
  wire  _GEN_395; // @[TLB.scala 251:68]
  wire  _GEN_396; // @[TLB.scala 251:68]
  wire  _GEN_403; // @[TLB.scala 251:68]
  wire  _GEN_404; // @[TLB.scala 251:68]
  wire  _GEN_405; // @[TLB.scala 251:68]
  wire  _GEN_406; // @[TLB.scala 251:68]
  wire  _GEN_413; // @[TLB.scala 251:68]
  wire  _GEN_414; // @[TLB.scala 251:68]
  wire  _GEN_415; // @[TLB.scala 251:68]
  wire  _GEN_416; // @[TLB.scala 251:68]
  wire  _GEN_423; // @[TLB.scala 251:68]
  wire  _GEN_424; // @[TLB.scala 251:68]
  wire  _GEN_425; // @[TLB.scala 251:68]
  wire  _GEN_426; // @[TLB.scala 251:68]
  wire  _GEN_433; // @[TLB.scala 251:68]
  wire  _GEN_434; // @[TLB.scala 251:68]
  wire  _GEN_435; // @[TLB.scala 251:68]
  wire  _GEN_436; // @[TLB.scala 251:68]
  wire  _GEN_443; // @[TLB.scala 251:68]
  wire  _GEN_444; // @[TLB.scala 251:68]
  wire  _GEN_445; // @[TLB.scala 251:68]
  wire  _GEN_446; // @[TLB.scala 251:68]
  wire  _GEN_455; // @[TLB.scala 224:40]
  wire  _GEN_459; // @[TLB.scala 224:40]
  wire  _GEN_463; // @[TLB.scala 224:40]
  wire  _GEN_467; // @[TLB.scala 224:40]
  wire  _GEN_471; // @[TLB.scala 224:40]
  wire  _GEN_473; // @[TLB.scala 224:40]
  wire  _GEN_474; // @[TLB.scala 224:40]
  wire  _GEN_475; // @[TLB.scala 224:40]
  wire  _GEN_476; // @[TLB.scala 224:40]
  wire  _GEN_483; // @[TLB.scala 224:40]
  wire  _GEN_484; // @[TLB.scala 224:40]
  wire  _GEN_485; // @[TLB.scala 224:40]
  wire  _GEN_486; // @[TLB.scala 224:40]
  wire  _GEN_493; // @[TLB.scala 224:40]
  wire  _GEN_494; // @[TLB.scala 224:40]
  wire  _GEN_495; // @[TLB.scala 224:40]
  wire  _GEN_496; // @[TLB.scala 224:40]
  wire  _GEN_503; // @[TLB.scala 224:40]
  wire  _GEN_504; // @[TLB.scala 224:40]
  wire  _GEN_505; // @[TLB.scala 224:40]
  wire  _GEN_506; // @[TLB.scala 224:40]
  wire  _GEN_513; // @[TLB.scala 224:40]
  wire  _GEN_514; // @[TLB.scala 224:40]
  wire  _GEN_515; // @[TLB.scala 224:40]
  wire  _GEN_516; // @[TLB.scala 224:40]
  wire  _GEN_523; // @[TLB.scala 224:40]
  wire  _GEN_524; // @[TLB.scala 224:40]
  wire  _GEN_525; // @[TLB.scala 224:40]
  wire  _GEN_526; // @[TLB.scala 224:40]
  wire  _GEN_533; // @[TLB.scala 224:40]
  wire  _GEN_534; // @[TLB.scala 224:40]
  wire  _GEN_535; // @[TLB.scala 224:40]
  wire  _GEN_536; // @[TLB.scala 224:40]
  wire  _GEN_543; // @[TLB.scala 224:40]
  wire  _GEN_544; // @[TLB.scala 224:40]
  wire  _GEN_545; // @[TLB.scala 224:40]
  wire  _GEN_546; // @[TLB.scala 224:40]
  wire [5:0] _T_2136; // @[Cat.scala 30:58]
  wire [13:0] ptw_ae_array; // @[Cat.scala 30:58]
  wire [5:0] _T_2150; // @[Cat.scala 30:58]
  wire [12:0] _T_2157; // @[Cat.scala 30:58]
  wire [12:0] priv_x_ok; // @[TLB.scala 307:22]
  wire [5:0] _T_2214; // @[Cat.scala 30:58]
  wire [12:0] _T_2221; // @[Cat.scala 30:58]
  wire [12:0] _T_2250; // @[TLB.scala 310:39]
  wire [13:0] x_array; // @[Cat.scala 30:58]
  wire [1:0] _T_2280; // @[Bitwise.scala 72:12]
  wire [5:0] _T_2285; // @[Cat.scala 30:58]
  wire [13:0] _T_2292; // @[Cat.scala 30:58]
  wire [13:0] px_array; // @[TLB.scala 313:87]
  wire [1:0] _T_2333; // @[Bitwise.scala 72:12]
  wire [5:0] _T_2338; // @[Cat.scala 30:58]
  wire [13:0] c_array; // @[Cat.scala 30:58]
  wire  _T_2364; // @[TLB.scala 323:37]
  wire [26:0] _T_2365; // @[TLB.scala 323:53]
  wire  _T_2366; // @[TLB.scala 323:60]
  wire  _T_2367; // @[TLB.scala 323:44]
  wire  bad_va; // @[TLB.scala 321:27]
  wire [13:0] _T_2549; // @[TLB.scala 338:33]
  wire [13:0] pf_inst_array; // @[TLB.scala 338:23]
  wire  tlb_hit; // @[TLB.scala 340:27]
  wire  _T_2551; // @[TLB.scala 341:29]
  wire  tlb_miss; // @[TLB.scala 341:40]
  reg [6:0] _T_2554; // @[Replacement.scala 41:30]
  reg [31:0] _RAND_100;
  reg [2:0] _T_2556; // @[Replacement.scala 41:30]
  reg [31:0] _RAND_101;
  wire  _T_2557; // @[TLB.scala 345:22]
  wire  _T_2558; // @[package.scala 63:59]
  wire  _T_2559; // @[package.scala 63:59]
  wire  _T_2560; // @[package.scala 63:59]
  wire  _T_2561; // @[package.scala 63:59]
  wire  _T_2562; // @[package.scala 63:59]
  wire  _T_2563; // @[package.scala 63:59]
  wire  _T_2564; // @[package.scala 63:59]
  wire [7:0] _T_2571; // @[Cat.scala 30:58]
  wire  _T_2574; // @[OneHot.scala 28:14]
  wire [3:0] _T_2575; // @[OneHot.scala 28:28]
  wire  _T_2578; // @[OneHot.scala 28:14]
  wire [1:0] _T_2579; // @[OneHot.scala 28:28]
  wire [2:0] _T_2582; // @[Cat.scala 30:58]
  wire [7:0] _T_2583; // @[Replacement.scala 46:28]
  wire [7:0] _T_2587; // @[Replacement.scala 50:37]
  wire [7:0] _T_2589; // @[Replacement.scala 50:37]
  wire [7:0] _T_2591; // @[Replacement.scala 50:37]
  wire [1:0] _T_2592; // @[Cat.scala 30:58]
  wire [3:0] _T_2595; // @[Replacement.scala 50:37]
  wire [7:0] _GEN_1001; // @[Replacement.scala 50:37]
  wire [7:0] _T_2596; // @[Replacement.scala 50:37]
  wire [7:0] _T_2598; // @[Replacement.scala 50:37]
  wire [7:0] _T_2600; // @[Replacement.scala 50:37]
  wire [2:0] _T_2601; // @[Cat.scala 30:58]
  wire [7:0] _T_2604; // @[Replacement.scala 50:37]
  wire [7:0] _T_2605; // @[Replacement.scala 50:37]
  wire [7:0] _T_2607; // @[Replacement.scala 50:37]
  wire [7:0] _T_2609; // @[Replacement.scala 50:37]
  wire  _T_2612; // @[package.scala 63:59]
  wire  _T_2613; // @[package.scala 63:59]
  wire  _T_2614; // @[package.scala 63:59]
  wire [3:0] _T_2617; // @[Cat.scala 30:58]
  wire  _T_2620; // @[OneHot.scala 28:14]
  wire [1:0] _T_2621; // @[OneHot.scala 28:28]
  wire [1:0] _T_2623; // @[Cat.scala 30:58]
  wire [3:0] _T_2624; // @[Replacement.scala 46:28]
  wire [3:0] _T_2628; // @[Replacement.scala 50:37]
  wire [3:0] _T_2630; // @[Replacement.scala 50:37]
  wire [3:0] _T_2632; // @[Replacement.scala 50:37]
  wire [1:0] _T_2633; // @[Cat.scala 30:58]
  wire [3:0] _T_2636; // @[Replacement.scala 50:37]
  wire [3:0] _T_2637; // @[Replacement.scala 50:37]
  wire [3:0] _T_2639; // @[Replacement.scala 50:37]
  wire [3:0] _T_2641; // @[Replacement.scala 50:37]
  wire  _T_2653; // @[Misc.scala 187:16]
  wire  _T_2655; // @[Misc.scala 187:61]
  wire  _T_2657; // @[Misc.scala 187:16]
  wire  _T_2659; // @[Misc.scala 187:61]
  wire  _T_2660; // @[Misc.scala 187:49]
  wire  _T_2669; // @[Misc.scala 187:16]
  wire  _T_2671; // @[Misc.scala 187:61]
  wire  _T_2673; // @[Misc.scala 187:16]
  wire  _T_2675; // @[Misc.scala 187:61]
  wire  _T_2676; // @[Misc.scala 187:49]
  wire  _T_2677; // @[Misc.scala 187:16]
  wire  _T_2678; // @[Misc.scala 187:37]
  wire  _T_2679; // @[Misc.scala 187:61]
  wire  _T_2680; // @[Misc.scala 187:49]
  wire  _T_2690; // @[Misc.scala 187:16]
  wire  _T_2692; // @[Misc.scala 187:61]
  wire  _T_2694; // @[Misc.scala 187:16]
  wire  _T_2696; // @[Misc.scala 187:61]
  wire  _T_2697; // @[Misc.scala 187:49]
  wire  _T_2704; // @[Misc.scala 187:16]
  wire  _T_2706; // @[Misc.scala 187:61]
  wire  _T_2713; // @[Misc.scala 187:16]
  wire  _T_2715; // @[Misc.scala 187:61]
  wire  _T_2717; // @[Misc.scala 187:16]
  wire  _T_2718; // @[Misc.scala 187:37]
  wire  _T_2719; // @[Misc.scala 187:61]
  wire  _T_2720; // @[Misc.scala 187:49]
  wire  _T_2721; // @[Misc.scala 187:16]
  wire  _T_2722; // @[Misc.scala 187:37]
  wire  _T_2723; // @[Misc.scala 187:61]
  wire  _T_2724; // @[Misc.scala 187:49]
  wire  _T_2726; // @[Misc.scala 187:37]
  wire  _T_2727; // @[Misc.scala 187:61]
  wire  multipleHits; // @[Misc.scala 187:49]
  wire [13:0] _T_2783; // @[TLB.scala 360:47]
  wire  _T_2784; // @[TLB.scala 360:55]
  wire [13:0] _T_2791; // @[TLB.scala 363:33]
  wire [13:0] _T_2797; // @[TLB.scala 367:33]
  wire  _T_2802; // @[TLB.scala 369:29]
  wire  _T_2808; // @[Decoupled.scala 37:37]
  wire  _T_2809; // @[TLB.scala 385:25]
  wire [3:0] _T_2814; // @[Replacement.scala 61:48]
  wire [1:0] _T_2817; // @[Cat.scala 30:58]
  wire [3:0] _T_2821; // @[Replacement.scala 61:48]
  wire [2:0] _T_2824; // @[Cat.scala 30:58]
  wire [3:0] _T_2828; // @[Cat.scala 30:58]
  wire  _T_2830; // @[TLB.scala 440:16]
  wire  _T_2832; // @[OneHot.scala 39:40]
  wire  _T_2833; // @[OneHot.scala 39:40]
  wire  _T_2834; // @[OneHot.scala 39:40]
  wire [7:0] _T_2844; // @[Replacement.scala 61:48]
  wire [1:0] _T_2847; // @[Cat.scala 30:58]
  wire [7:0] _T_2851; // @[Replacement.scala 61:48]
  wire [2:0] _T_2854; // @[Cat.scala 30:58]
  wire [7:0] _T_2858; // @[Replacement.scala 61:48]
  wire [3:0] _T_2861; // @[Cat.scala 30:58]
  wire [7:0] _T_2893; // @[Cat.scala 30:58]
  wire  _T_2895; // @[TLB.scala 440:16]
  wire  _T_2897; // @[OneHot.scala 39:40]
  wire  _T_2898; // @[OneHot.scala 39:40]
  wire  _T_2899; // @[OneHot.scala 39:40]
  wire  _T_2900; // @[OneHot.scala 39:40]
  wire  _T_2901; // @[OneHot.scala 39:40]
  wire  _T_2902; // @[OneHot.scala 39:40]
  wire  _T_2903; // @[OneHot.scala 39:40]
  wire  _T_2940; // @[TLB.scala 399:17]
  wire  _T_2941; // @[TLB.scala 399:28]
  wire  _T_2946; // @[TLB.scala 414:72]
  wire  _T_2947; // @[TLB.scala 414:34]
  wire  _T_2949; // @[TLB.scala 414:13]
  wire  _T_2957; // @[TLB.scala 150:63]
  wire  _GEN_652; // @[TLB.scala 158:21]
  wire  _GEN_653; // @[TLB.scala 158:21]
  wire  _GEN_654; // @[TLB.scala 158:21]
  wire  _GEN_655; // @[TLB.scala 158:21]
  wire  _GEN_656; // @[TLB.scala 417:40]
  wire  _GEN_657; // @[TLB.scala 417:40]
  wire  _GEN_658; // @[TLB.scala 417:40]
  wire  _GEN_659; // @[TLB.scala 417:40]
  wire  _T_3128; // @[TLB.scala 150:63]
  wire  _GEN_680; // @[TLB.scala 158:21]
  wire  _GEN_681; // @[TLB.scala 158:21]
  wire  _GEN_682; // @[TLB.scala 158:21]
  wire  _GEN_683; // @[TLB.scala 158:21]
  wire  _GEN_684; // @[TLB.scala 417:40]
  wire  _GEN_685; // @[TLB.scala 417:40]
  wire  _GEN_686; // @[TLB.scala 417:40]
  wire  _GEN_687; // @[TLB.scala 417:40]
  wire  _T_3299; // @[TLB.scala 150:63]
  wire  _GEN_708; // @[TLB.scala 158:21]
  wire  _GEN_709; // @[TLB.scala 158:21]
  wire  _GEN_710; // @[TLB.scala 158:21]
  wire  _GEN_711; // @[TLB.scala 158:21]
  wire  _GEN_712; // @[TLB.scala 417:40]
  wire  _GEN_713; // @[TLB.scala 417:40]
  wire  _GEN_714; // @[TLB.scala 417:40]
  wire  _GEN_715; // @[TLB.scala 417:40]
  wire  _T_3470; // @[TLB.scala 150:63]
  wire  _GEN_736; // @[TLB.scala 158:21]
  wire  _GEN_737; // @[TLB.scala 158:21]
  wire  _GEN_738; // @[TLB.scala 158:21]
  wire  _GEN_739; // @[TLB.scala 158:21]
  wire  _GEN_740; // @[TLB.scala 417:40]
  wire  _GEN_741; // @[TLB.scala 417:40]
  wire  _GEN_742; // @[TLB.scala 417:40]
  wire  _GEN_743; // @[TLB.scala 417:40]
  wire  _T_3641; // @[TLB.scala 150:63]
  wire  _GEN_764; // @[TLB.scala 158:21]
  wire  _GEN_765; // @[TLB.scala 158:21]
  wire  _GEN_766; // @[TLB.scala 158:21]
  wire  _GEN_767; // @[TLB.scala 158:21]
  wire  _GEN_768; // @[TLB.scala 417:40]
  wire  _GEN_769; // @[TLB.scala 417:40]
  wire  _GEN_770; // @[TLB.scala 417:40]
  wire  _GEN_771; // @[TLB.scala 417:40]
  wire  _T_3812; // @[TLB.scala 150:63]
  wire  _GEN_792; // @[TLB.scala 158:21]
  wire  _GEN_793; // @[TLB.scala 158:21]
  wire  _GEN_794; // @[TLB.scala 158:21]
  wire  _GEN_795; // @[TLB.scala 158:21]
  wire  _GEN_796; // @[TLB.scala 417:40]
  wire  _GEN_797; // @[TLB.scala 417:40]
  wire  _GEN_798; // @[TLB.scala 417:40]
  wire  _GEN_799; // @[TLB.scala 417:40]
  wire  _T_3983; // @[TLB.scala 150:63]
  wire  _GEN_820; // @[TLB.scala 158:21]
  wire  _GEN_821; // @[TLB.scala 158:21]
  wire  _GEN_822; // @[TLB.scala 158:21]
  wire  _GEN_823; // @[TLB.scala 158:21]
  wire  _GEN_824; // @[TLB.scala 417:40]
  wire  _GEN_825; // @[TLB.scala 417:40]
  wire  _GEN_826; // @[TLB.scala 417:40]
  wire  _GEN_827; // @[TLB.scala 417:40]
  wire  _T_4154; // @[TLB.scala 150:63]
  wire  _GEN_848; // @[TLB.scala 158:21]
  wire  _GEN_849; // @[TLB.scala 158:21]
  wire  _GEN_850; // @[TLB.scala 158:21]
  wire  _GEN_851; // @[TLB.scala 158:21]
  wire  _GEN_852; // @[TLB.scala 417:40]
  wire  _GEN_853; // @[TLB.scala 417:40]
  wire  _GEN_854; // @[TLB.scala 417:40]
  wire  _GEN_855; // @[TLB.scala 417:40]
  wire  _GEN_861; // @[TLB.scala 158:21]
  wire  _GEN_862; // @[TLB.scala 417:40]
  wire  _GEN_865; // @[TLB.scala 158:21]
  wire  _GEN_866; // @[TLB.scala 417:40]
  wire  _GEN_869; // @[TLB.scala 158:21]
  wire  _GEN_870; // @[TLB.scala 417:40]
  wire  _GEN_873; // @[TLB.scala 158:21]
  wire  _GEN_874; // @[TLB.scala 417:40]
  wire  _GEN_877; // @[TLB.scala 158:21]
  wire  _GEN_878; // @[TLB.scala 417:40]
  wire  _T_4530; // @[TLB.scala 421:24]
  reg [19:0] TLB_1_state; // @[Register tracking TLB_1 state]
  reg [31:0] _RAND_102;
  reg  TLB_1_cov [0:1048575]; // @[Coverage map for TLB_1]
  reg [31:0] _RAND_103;
  wire  TLB_1_cov_read_data; // @[Coverage map for TLB_1]
  wire [19:0] TLB_1_cov_read_addr; // @[Coverage map for TLB_1]
  wire  TLB_1_cov_write_data; // @[Coverage map for TLB_1]
  wire [19:0] TLB_1_cov_write_addr; // @[Coverage map for TLB_1]
  wire  TLB_1_cov_write_mask; // @[Coverage map for TLB_1]
  wire  TLB_1_cov_write_en; // @[Coverage map for TLB_1]
  reg [29:0] TLB_1_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_104;
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  mux_cond_4;
  wire  mux_cond_5;
  wire  mux_cond_6;
  wire  mux_cond_7;
  wire  mux_cond_8;
  wire  mux_cond_9;
  wire  mux_cond_10;
  wire  mux_cond_11;
  wire  mux_cond_12;
  wire  mux_cond_13;
  wire  mux_cond_14;
  wire  mux_cond_15;
  wire  mux_cond_16;
  wire  mux_cond_17;
  wire  mux_cond_18;
  wire  mux_cond_19;
  wire  mux_cond_20;
  wire  mux_cond_21;
  wire  mux_cond_22;
  wire  mux_cond_23;
  wire  mux_cond_24;
  wire  mux_cond_25;
  wire  mux_cond_26;
  wire  mux_cond_27;
  wire  mux_cond_28;
  wire  mux_cond_29;
  wire  mux_cond_30;
  wire  mux_cond_31;
  wire  mux_cond_32;
  wire  mux_cond_33;
  wire  mux_cond_34;
  wire  mux_cond_35;
  wire  mux_cond_36;
  wire  mux_cond_37;
  wire  mux_cond_38;
  wire  mux_cond_39;
  wire  mux_cond_40;
  wire  mux_cond_41;
  wire  mux_cond_42;
  wire  mux_cond_43;
  wire  mux_cond_44;
  wire  mux_cond_45;
  wire  mux_cond_46;
  wire  mux_cond_47;
  wire  mux_cond_48;
  wire  mux_cond_49;
  wire  mux_cond_50;
  wire  mux_cond_51;
  wire  mux_cond_52;
  wire  mux_cond_53;
  wire  mux_cond_54;
  wire  mux_cond_55;
  wire  mux_cond_56;
  wire  mux_cond_57;
  wire  mux_cond_58;
  wire  mux_cond_59;
  wire  mux_cond_60;
  wire  mux_cond_61;
  wire  mux_cond_62;
  wire  mux_cond_63;
  wire  mux_cond_64;
  wire  mux_cond_65;
  wire  mux_cond_66;
  wire  mux_cond_67;
  wire  mux_cond_68;
  wire  mux_cond_69;
  wire  mux_cond_70;
  wire [19:0] r_superpage_repl_addr_shl;
  wire [19:0] r_superpage_repl_addr_pad;
  wire [4:0] state_shl;
  wire [19:0] state_pad;
  wire [16:0] r_sectored_repl_addr_shl;
  wire [19:0] r_sectored_repl_addr_pad;
  wire [5:0] r_sectored_hit_addr_shl;
  wire [19:0] r_sectored_hit_addr_pad;
  wire [9:0] special_entry_valid_0_shl;
  wire [19:0] special_entry_valid_0_pad;
  wire [2:0] special_entry_level_shl;
  wire [19:0] special_entry_level_pad;
  wire [1:0] r_sectored_hit_shl;
  wire [19:0] r_sectored_hit_pad;
  wire [1:0] mux_cond_0_shl;
  wire [19:0] mux_cond_0_pad;
  wire [3:0] mux_cond_1_shl;
  wire [19:0] mux_cond_1_pad;
  wire [6:0] mux_cond_2_shl;
  wire [19:0] mux_cond_2_pad;
  wire [14:0] mux_cond_3_shl;
  wire [19:0] mux_cond_3_pad;
  wire [17:0] mux_cond_4_shl;
  wire [19:0] mux_cond_4_pad;
  wire [19:0] mux_cond_5_shl;
  wire [19:0] mux_cond_5_pad;
  wire [7:0] mux_cond_6_shl;
  wire [19:0] mux_cond_6_pad;
  wire [16:0] mux_cond_7_shl;
  wire [19:0] mux_cond_7_pad;
  wire [7:0] mux_cond_8_shl;
  wire [19:0] mux_cond_8_pad;
  wire [10:0] mux_cond_9_shl;
  wire [19:0] mux_cond_9_pad;
  wire [14:0] mux_cond_10_shl;
  wire [19:0] mux_cond_10_pad;
  wire [9:0] mux_cond_11_shl;
  wire [19:0] mux_cond_11_pad;
  wire [9:0] mux_cond_12_shl;
  wire [19:0] mux_cond_12_pad;
  wire [9:0] mux_cond_13_shl;
  wire [19:0] mux_cond_13_pad;
  wire [14:0] mux_cond_14_shl;
  wire [19:0] mux_cond_14_pad;
  wire [8:0] mux_cond_15_shl;
  wire [19:0] mux_cond_15_pad;
  wire [15:0] mux_cond_16_shl;
  wire [19:0] mux_cond_16_pad;
  wire [10:0] mux_cond_17_shl;
  wire [19:0] mux_cond_17_pad;
  wire  mux_cond_18_shl;
  wire [19:0] mux_cond_18_pad;
  wire [13:0] mux_cond_19_shl;
  wire [19:0] mux_cond_19_pad;
  wire [9:0] mux_cond_20_shl;
  wire [19:0] mux_cond_20_pad;
  wire [16:0] mux_cond_21_shl;
  wire [19:0] mux_cond_21_pad;
  wire [5:0] mux_cond_22_shl;
  wire [19:0] mux_cond_22_pad;
  wire [19:0] mux_cond_23_shl;
  wire [19:0] mux_cond_23_pad;
  wire [1:0] mux_cond_24_shl;
  wire [19:0] mux_cond_24_pad;
  wire [8:0] mux_cond_25_shl;
  wire [19:0] mux_cond_25_pad;
  wire [12:0] mux_cond_26_shl;
  wire [19:0] mux_cond_26_pad;
  wire [14:0] mux_cond_27_shl;
  wire [19:0] mux_cond_27_pad;
  wire [7:0] mux_cond_28_shl;
  wire [19:0] mux_cond_28_pad;
  wire [11:0] mux_cond_29_shl;
  wire [19:0] mux_cond_29_pad;
  wire [8:0] mux_cond_30_shl;
  wire [19:0] mux_cond_30_pad;
  wire [6:0] mux_cond_31_shl;
  wire [19:0] mux_cond_31_pad;
  wire [6:0] mux_cond_32_shl;
  wire [19:0] mux_cond_32_pad;
  wire [6:0] mux_cond_33_shl;
  wire [19:0] mux_cond_33_pad;
  wire [16:0] mux_cond_34_shl;
  wire [19:0] mux_cond_34_pad;
  wire [11:0] mux_cond_35_shl;
  wire [19:0] mux_cond_35_pad;
  wire [4:0] mux_cond_36_shl;
  wire [19:0] mux_cond_36_pad;
  wire [7:0] mux_cond_37_shl;
  wire [19:0] mux_cond_37_pad;
  wire [11:0] mux_cond_38_shl;
  wire [19:0] mux_cond_38_pad;
  wire [14:0] mux_cond_39_shl;
  wire [19:0] mux_cond_39_pad;
  wire [7:0] mux_cond_40_shl;
  wire [19:0] mux_cond_40_pad;
  wire [9:0] mux_cond_41_shl;
  wire [19:0] mux_cond_41_pad;
  wire [1:0] mux_cond_42_shl;
  wire [19:0] mux_cond_42_pad;
  wire [4:0] mux_cond_43_shl;
  wire [19:0] mux_cond_43_pad;
  wire [6:0] mux_cond_44_shl;
  wire [19:0] mux_cond_44_pad;
  wire [15:0] mux_cond_45_shl;
  wire [19:0] mux_cond_45_pad;
  wire [18:0] mux_cond_46_shl;
  wire [19:0] mux_cond_46_pad;
  wire [2:0] mux_cond_47_shl;
  wire [19:0] mux_cond_47_pad;
  wire [11:0] mux_cond_48_shl;
  wire [19:0] mux_cond_48_pad;
  wire [14:0] mux_cond_49_shl;
  wire [19:0] mux_cond_49_pad;
  wire [15:0] mux_cond_50_shl;
  wire [19:0] mux_cond_50_pad;
  wire [9:0] mux_cond_51_shl;
  wire [19:0] mux_cond_51_pad;
  wire [18:0] mux_cond_52_shl;
  wire [19:0] mux_cond_52_pad;
  wire [18:0] mux_cond_53_shl;
  wire [19:0] mux_cond_53_pad;
  wire [10:0] mux_cond_54_shl;
  wire [19:0] mux_cond_54_pad;
  wire [9:0] mux_cond_55_shl;
  wire [19:0] mux_cond_55_pad;
  wire  mux_cond_56_shl;
  wire [19:0] mux_cond_56_pad;
  wire [3:0] mux_cond_57_shl;
  wire [19:0] mux_cond_57_pad;
  wire [19:0] mux_cond_58_shl;
  wire [19:0] mux_cond_58_pad;
  wire [2:0] mux_cond_59_shl;
  wire [19:0] mux_cond_59_pad;
  wire [15:0] mux_cond_60_shl;
  wire [19:0] mux_cond_60_pad;
  wire [17:0] mux_cond_61_shl;
  wire [19:0] mux_cond_61_pad;
  wire [11:0] mux_cond_62_shl;
  wire [19:0] mux_cond_62_pad;
  wire [15:0] mux_cond_63_shl;
  wire [19:0] mux_cond_63_pad;
  wire [9:0] mux_cond_64_shl;
  wire [19:0] mux_cond_64_pad;
  wire [17:0] mux_cond_65_shl;
  wire [19:0] mux_cond_65_pad;
  wire [12:0] mux_cond_66_shl;
  wire [19:0] mux_cond_66_pad;
  wire [15:0] mux_cond_67_shl;
  wire [19:0] mux_cond_67_pad;
  wire [17:0] mux_cond_68_shl;
  wire [19:0] mux_cond_68_pad;
  wire [3:0] mux_cond_69_shl;
  wire [19:0] mux_cond_69_pad;
  wire [3:0] mux_cond_70_shl;
  wire [19:0] mux_cond_70_pad;
  wire [12:0] sectored_entries_7_valid_1_shl;
  wire [19:0] sectored_entries_7_valid_1_pad;
  wire [7:0] sectored_entries_5_valid_3_shl;
  wire [19:0] sectored_entries_5_valid_3_pad;
  wire [12:0] sectored_entries_5_valid_1_shl;
  wire [19:0] sectored_entries_5_valid_1_pad;
  wire [12:0] sectored_entries_4_valid_1_shl;
  wire [19:0] sectored_entries_4_valid_1_pad;
  wire [6:0] superpage_entries_0_valid_0_shl;
  wire [19:0] superpage_entries_0_valid_0_pad;
  wire [9:0] sectored_entries_3_valid_2_shl;
  wire [19:0] sectored_entries_3_valid_2_pad;
  wire [9:0] sectored_entries_1_valid_0_shl;
  wire [19:0] sectored_entries_1_valid_0_pad;
  wire [3:0] superpage_entries_3_level_shl;
  wire [19:0] superpage_entries_3_level_pad;
  wire [9:0] sectored_entries_5_valid_0_shl;
  wire [19:0] sectored_entries_5_valid_0_pad;
  wire [12:0] sectored_entries_0_valid_1_shl;
  wire [19:0] sectored_entries_0_valid_1_pad;
  wire [9:0] sectored_entries_3_valid_0_shl;
  wire [19:0] sectored_entries_3_valid_0_pad;
  wire [9:0] sectored_entries_7_valid_2_shl;
  wire [19:0] sectored_entries_7_valid_2_pad;
  wire [7:0] sectored_entries_2_valid_3_shl;
  wire [19:0] sectored_entries_2_valid_3_pad;
  wire [9:0] sectored_entries_4_valid_0_shl;
  wire [19:0] sectored_entries_4_valid_0_pad;
  wire [7:0] sectored_entries_6_valid_3_shl;
  wire [19:0] sectored_entries_6_valid_3_pad;
  wire [7:0] sectored_entries_1_valid_3_shl;
  wire [19:0] sectored_entries_1_valid_3_pad;
  wire [9:0] sectored_entries_6_valid_0_shl;
  wire [19:0] sectored_entries_6_valid_0_pad;
  wire [9:0] sectored_entries_2_valid_2_shl;
  wire [19:0] sectored_entries_2_valid_2_pad;
  wire [9:0] sectored_entries_6_valid_2_shl;
  wire [19:0] sectored_entries_6_valid_2_pad;
  wire [12:0] sectored_entries_6_valid_1_shl;
  wire [19:0] sectored_entries_6_valid_1_pad;
  wire [7:0] sectored_entries_4_valid_3_shl;
  wire [19:0] sectored_entries_4_valid_3_pad;
  wire [9:0] sectored_entries_1_valid_2_shl;
  wire [19:0] sectored_entries_1_valid_2_pad;
  wire [9:0] sectored_entries_5_valid_2_shl;
  wire [19:0] sectored_entries_5_valid_2_pad;
  wire [3:0] superpage_entries_2_level_shl;
  wire [19:0] superpage_entries_2_level_pad;
  wire [6:0] superpage_entries_3_valid_0_shl;
  wire [19:0] superpage_entries_3_valid_0_pad;
  wire [12:0] sectored_entries_1_valid_1_shl;
  wire [19:0] sectored_entries_1_valid_1_pad;
  wire [9:0] sectored_entries_0_valid_0_shl;
  wire [19:0] sectored_entries_0_valid_0_pad;
  wire [6:0] superpage_entries_1_valid_0_shl;
  wire [19:0] superpage_entries_1_valid_0_pad;
  wire [7:0] sectored_entries_0_valid_3_shl;
  wire [19:0] sectored_entries_0_valid_3_pad;
  wire [9:0] sectored_entries_7_valid_0_shl;
  wire [19:0] sectored_entries_7_valid_0_pad;
  wire [9:0] sectored_entries_0_valid_2_shl;
  wire [19:0] sectored_entries_0_valid_2_pad;
  wire [3:0] superpage_entries_0_level_shl;
  wire [19:0] superpage_entries_0_level_pad;
  wire [12:0] sectored_entries_2_valid_1_shl;
  wire [19:0] sectored_entries_2_valid_1_pad;
  wire [12:0] sectored_entries_3_valid_1_shl;
  wire [19:0] sectored_entries_3_valid_1_pad;
  wire [9:0] sectored_entries_2_valid_0_shl;
  wire [19:0] sectored_entries_2_valid_0_pad;
  wire [7:0] sectored_entries_7_valid_3_shl;
  wire [19:0] sectored_entries_7_valid_3_pad;
  wire [9:0] sectored_entries_4_valid_2_shl;
  wire [19:0] sectored_entries_4_valid_2_pad;
  wire [7:0] sectored_entries_3_valid_3_shl;
  wire [19:0] sectored_entries_3_valid_3_pad;
  wire [3:0] superpage_entries_1_level_shl;
  wire [19:0] superpage_entries_1_level_pad;
  wire [6:0] superpage_entries_2_valid_0_shl;
  wire [19:0] superpage_entries_2_valid_0_pad;
  wire [19:0] TLB_1_xor64;
  wire [19:0] TLB_1_xor31;
  wire [19:0] TLB_1_xor65;
  wire [19:0] TLB_1_xor66;
  wire [19:0] TLB_1_xor32;
  wire [19:0] TLB_1_xor15;
  wire [19:0] TLB_1_xor68;
  wire [19:0] TLB_1_xor33;
  wire [19:0] TLB_1_xor69;
  wire [19:0] TLB_1_xor70;
  wire [19:0] TLB_1_xor34;
  wire [19:0] TLB_1_xor16;
  wire [19:0] TLB_1_xor7;
  wire [19:0] TLB_1_xor72;
  wire [19:0] TLB_1_xor35;
  wire [19:0] TLB_1_xor73;
  wire [19:0] TLB_1_xor74;
  wire [19:0] TLB_1_xor36;
  wire [19:0] TLB_1_xor17;
  wire [19:0] TLB_1_xor75;
  wire [19:0] TLB_1_xor76;
  wire [19:0] TLB_1_xor37;
  wire [19:0] TLB_1_xor77;
  wire [19:0] TLB_1_xor78;
  wire [19:0] TLB_1_xor38;
  wire [19:0] TLB_1_xor18;
  wire [19:0] TLB_1_xor8;
  wire [19:0] TLB_1_xor3;
  wire [19:0] TLB_1_xor80;
  wire [19:0] TLB_1_xor39;
  wire [19:0] TLB_1_xor81;
  wire [19:0] TLB_1_xor82;
  wire [19:0] TLB_1_xor40;
  wire [19:0] TLB_1_xor19;
  wire [19:0] TLB_1_xor83;
  wire [19:0] TLB_1_xor84;
  wire [19:0] TLB_1_xor41;
  wire [19:0] TLB_1_xor85;
  wire [19:0] TLB_1_xor86;
  wire [19:0] TLB_1_xor42;
  wire [19:0] TLB_1_xor20;
  wire [19:0] TLB_1_xor9;
  wire [19:0] TLB_1_xor88;
  wire [19:0] TLB_1_xor43;
  wire [19:0] TLB_1_xor89;
  wire [19:0] TLB_1_xor90;
  wire [19:0] TLB_1_xor44;
  wire [19:0] TLB_1_xor21;
  wire [19:0] TLB_1_xor91;
  wire [19:0] TLB_1_xor92;
  wire [19:0] TLB_1_xor45;
  wire [19:0] TLB_1_xor93;
  wire [19:0] TLB_1_xor94;
  wire [19:0] TLB_1_xor46;
  wire [19:0] TLB_1_xor22;
  wire [19:0] TLB_1_xor10;
  wire [19:0] TLB_1_xor4;
  wire [19:0] TLB_1_xor1;
  wire [19:0] TLB_1_xor96;
  wire [19:0] TLB_1_xor47;
  wire [19:0] TLB_1_xor97;
  wire [19:0] TLB_1_xor98;
  wire [19:0] TLB_1_xor48;
  wire [19:0] TLB_1_xor23;
  wire [19:0] TLB_1_xor100;
  wire [19:0] TLB_1_xor49;
  wire [19:0] TLB_1_xor101;
  wire [19:0] TLB_1_xor102;
  wire [19:0] TLB_1_xor50;
  wire [19:0] TLB_1_xor24;
  wire [19:0] TLB_1_xor11;
  wire [19:0] TLB_1_xor104;
  wire [19:0] TLB_1_xor51;
  wire [19:0] TLB_1_xor105;
  wire [19:0] TLB_1_xor106;
  wire [19:0] TLB_1_xor52;
  wire [19:0] TLB_1_xor25;
  wire [19:0] TLB_1_xor107;
  wire [19:0] TLB_1_xor108;
  wire [19:0] TLB_1_xor53;
  wire [19:0] TLB_1_xor109;
  wire [19:0] TLB_1_xor110;
  wire [19:0] TLB_1_xor54;
  wire [19:0] TLB_1_xor26;
  wire [19:0] TLB_1_xor12;
  wire [19:0] TLB_1_xor5;
  wire [19:0] TLB_1_xor112;
  wire [19:0] TLB_1_xor55;
  wire [19:0] TLB_1_xor113;
  wire [19:0] TLB_1_xor114;
  wire [19:0] TLB_1_xor56;
  wire [19:0] TLB_1_xor27;
  wire [19:0] TLB_1_xor115;
  wire [19:0] TLB_1_xor116;
  wire [19:0] TLB_1_xor57;
  wire [19:0] TLB_1_xor117;
  wire [19:0] TLB_1_xor118;
  wire [19:0] TLB_1_xor58;
  wire [19:0] TLB_1_xor28;
  wire [19:0] TLB_1_xor13;
  wire [19:0] TLB_1_xor120;
  wire [19:0] TLB_1_xor59;
  wire [19:0] TLB_1_xor121;
  wire [19:0] TLB_1_xor122;
  wire [19:0] TLB_1_xor60;
  wire [19:0] TLB_1_xor29;
  wire [19:0] TLB_1_xor123;
  wire [19:0] TLB_1_xor124;
  wire [19:0] TLB_1_xor61;
  wire [19:0] TLB_1_xor125;
  wire [19:0] TLB_1_xor126;
  wire [19:0] TLB_1_xor62;
  wire [19:0] TLB_1_xor30;
  wire [19:0] TLB_1_xor14;
  wire [19:0] TLB_1_xor6;
  wire [19:0] TLB_1_xor2;
  wire [19:0] TLB_1_xor0;
  wire [29:0] pmp_sum;
  wire  stopEn0;
  wire  pmp_metaAssert_wire;
  wire  TLB_1_or0;
  reg  TLB_1_metaAssert;
  reg [31:0] _RAND_105;
  PMPChecker_1 pmp ( // @[TLB.scala 190:19]
    .io_prv(pmp_io_prv),
    .io_pmp_0_cfg_l(pmp_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(pmp_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(pmp_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(pmp_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(pmp_io_pmp_0_cfg_r),
    .io_pmp_0_addr(pmp_io_pmp_0_addr),
    .io_pmp_0_mask(pmp_io_pmp_0_mask),
    .io_pmp_1_cfg_l(pmp_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(pmp_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(pmp_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(pmp_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(pmp_io_pmp_1_cfg_r),
    .io_pmp_1_addr(pmp_io_pmp_1_addr),
    .io_pmp_1_mask(pmp_io_pmp_1_mask),
    .io_pmp_2_cfg_l(pmp_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(pmp_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(pmp_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(pmp_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(pmp_io_pmp_2_cfg_r),
    .io_pmp_2_addr(pmp_io_pmp_2_addr),
    .io_pmp_2_mask(pmp_io_pmp_2_mask),
    .io_pmp_3_cfg_l(pmp_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(pmp_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(pmp_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(pmp_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(pmp_io_pmp_3_cfg_r),
    .io_pmp_3_addr(pmp_io_pmp_3_addr),
    .io_pmp_3_mask(pmp_io_pmp_3_mask),
    .io_pmp_4_cfg_l(pmp_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(pmp_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(pmp_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(pmp_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(pmp_io_pmp_4_cfg_r),
    .io_pmp_4_addr(pmp_io_pmp_4_addr),
    .io_pmp_4_mask(pmp_io_pmp_4_mask),
    .io_pmp_5_cfg_l(pmp_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(pmp_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(pmp_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(pmp_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(pmp_io_pmp_5_cfg_r),
    .io_pmp_5_addr(pmp_io_pmp_5_addr),
    .io_pmp_5_mask(pmp_io_pmp_5_mask),
    .io_pmp_6_cfg_l(pmp_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(pmp_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(pmp_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(pmp_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(pmp_io_pmp_6_cfg_r),
    .io_pmp_6_addr(pmp_io_pmp_6_addr),
    .io_pmp_6_mask(pmp_io_pmp_6_mask),
    .io_pmp_7_cfg_l(pmp_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(pmp_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(pmp_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(pmp_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(pmp_io_pmp_7_cfg_r),
    .io_pmp_7_addr(pmp_io_pmp_7_addr),
    .io_pmp_7_mask(pmp_io_pmp_7_mask),
    .io_addr(pmp_io_addr),
    .io_r(pmp_io_r),
    .io_w(pmp_io_w),
    .io_x(pmp_io_x),
    .io_covSum(pmp_io_covSum),
    .metaAssert(pmp_metaAssert)
  );
  assign priv_s = io_ptw_status_prv[0]; // @[TLB.scala 178:20]
  assign priv_uses_vm = io_ptw_status_prv <= 2'h1; // @[TLB.scala 179:27]
  assign vm_enabled = io_ptw_ptbr_mode[3] & priv_uses_vm; // @[TLB.scala 180:83]
  assign vpn = io_req_bits_vaddr[38:12]; // @[TLB.scala 183:30]
  assign refill_ppn = io_ptw_resp_bits_pte_ppn[19:0]; // @[TLB.scala 184:44]
  assign _T_324 = state == 2'h1; // @[package.scala 14:47]
  assign _T_325 = state == 2'h3; // @[package.scala 14:47]
  assign invalidate_refill = _T_324 | _T_325; // @[package.scala 14:62]
  assign _T_348 = special_entry_level < 2'h1; // @[TLB.scala 123:30]
  assign _T_350 = _T_348 ? vpn : 27'h0; // @[TLB.scala 124:30]
  assign _GEN_954 = {{7'd0}, special_entry_data_0[33:14]}; // @[TLB.scala 124:49]
  assign _T_351 = _T_350 | _GEN_954; // @[TLB.scala 124:49]
  assign _T_354 = special_entry_level < 2'h2; // @[TLB.scala 123:30]
  assign _T_356 = _T_354 ? vpn : 27'h0; // @[TLB.scala 124:30]
  assign _T_357 = _T_356 | _GEN_954; // @[TLB.scala 124:49]
  assign _T_359 = {special_entry_data_0[33:32],_T_351[17:9],_T_357[8:0]}; // @[Cat.scala 30:58]
  assign _T_361 = vm_enabled ? {{8'd0}, _T_359} : io_req_bits_vaddr[39:12]; // @[TLB.scala 188:20]
  assign mpu_ppn = io_ptw_resp_valid ? {{8'd0}, refill_ppn} : _T_361; // @[TLB.scala 187:20]
  assign mpu_physaddr = {mpu_ppn,io_req_bits_vaddr[11:0]}; // @[Cat.scala 30:58]
  assign _T_366 = mpu_physaddr ^ 40'h3000; // @[Parameters.scala 121:31]
  assign _T_367 = {1'b0,$signed(_T_366)}; // @[Parameters.scala 121:49]
  assign _T_369 = $signed(_T_367) & -41'sh1000; // @[Parameters.scala 121:52]
  assign _T_370 = $signed(_T_369) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_371 = mpu_physaddr ^ 40'hc000000; // @[Parameters.scala 121:31]
  assign _T_372 = {1'b0,$signed(_T_371)}; // @[Parameters.scala 121:49]
  assign _T_374 = $signed(_T_372) & -41'sh4000000; // @[Parameters.scala 121:52]
  assign _T_375 = $signed(_T_374) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_376 = mpu_physaddr ^ 40'h2000000; // @[Parameters.scala 121:31]
  assign _T_377 = {1'b0,$signed(_T_376)}; // @[Parameters.scala 121:49]
  assign _T_379 = $signed(_T_377) & -41'sh10000; // @[Parameters.scala 121:52]
  assign _T_380 = $signed(_T_379) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_382 = {1'b0,$signed(mpu_physaddr)}; // @[Parameters.scala 121:49]
  assign _T_384 = $signed(_T_382) & -41'sh1000; // @[Parameters.scala 121:52]
  assign _T_385 = $signed(_T_384) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_386 = mpu_physaddr ^ 40'h10000; // @[Parameters.scala 121:31]
  assign _T_387 = {1'b0,$signed(_T_386)}; // @[Parameters.scala 121:49]
  assign _T_389 = $signed(_T_387) & -41'sh10000; // @[Parameters.scala 121:52]
  assign _T_390 = $signed(_T_389) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_391 = mpu_physaddr ^ 40'h80000000; // @[Parameters.scala 121:31]
  assign _T_392 = {1'b0,$signed(_T_391)}; // @[Parameters.scala 121:49]
  assign _T_394 = $signed(_T_392) & -41'sh10000000; // @[Parameters.scala 121:52]
  assign _T_395 = $signed(_T_394) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_396 = mpu_physaddr ^ 40'h60000000; // @[Parameters.scala 121:31]
  assign _T_397 = {1'b0,$signed(_T_396)}; // @[Parameters.scala 121:49]
  assign _T_399 = $signed(_T_397) & -41'sh20000000; // @[Parameters.scala 121:52]
  assign _T_400 = $signed(_T_399) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_414 = _T_370 | _T_375; // @[TLB.scala 195:67]
  assign _T_415 = _T_414 | _T_380; // @[TLB.scala 195:67]
  assign _T_416 = _T_415 | _T_385; // @[TLB.scala 195:67]
  assign _T_417 = _T_416 | _T_390; // @[TLB.scala 195:67]
  assign _T_418 = _T_417 | _T_395; // @[TLB.scala 195:67]
  assign legal_address = _T_418 | _T_400; // @[TLB.scala 195:67]
  assign _T_427 = $signed(_T_392) & 41'sh80000000; // @[Parameters.scala 121:52]
  assign _T_428 = $signed(_T_427) == 41'sh0; // @[Parameters.scala 121:67]
  assign cacheable = legal_address & _T_428; // @[TLB.scala 197:19]
  assign _T_485 = mpu_physaddr ^ 40'h8000000; // @[Parameters.scala 121:31]
  assign _T_486 = {1'b0,$signed(_T_485)}; // @[Parameters.scala 121:49]
  assign _T_488 = $signed(_T_486) & 41'shc8000000; // @[Parameters.scala 121:52]
  assign _T_489 = $signed(_T_488) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_507 = $signed(_T_382) & 41'shc8010000; // @[Parameters.scala 121:52]
  assign _T_508 = $signed(_T_507) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_515 = _T_508 | _T_489; // @[TLBPermissions.scala 81:66]
  assign prot_r = legal_address & pmp_io_r; // @[TLB.scala 200:41]
  assign _T_552 = $signed(_T_392) & 41'shc0000000; // @[Parameters.scala 121:52]
  assign _T_553 = $signed(_T_552) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_554 = mpu_physaddr ^ 40'h40000000; // @[Parameters.scala 121:31]
  assign _T_555 = {1'b0,$signed(_T_554)}; // @[Parameters.scala 121:49]
  assign _T_557 = $signed(_T_555) & 41'shc0000000; // @[Parameters.scala 121:52]
  assign _T_558 = $signed(_T_557) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_560 = _T_515 | _T_553; // @[Parameters.scala 148:89]
  assign _T_561 = _T_560 | _T_558; // @[Parameters.scala 148:89]
  assign _T_568 = legal_address & _T_561; // @[TLB.scala 197:19]
  assign prot_w = _T_568 & pmp_io_w; // @[TLB.scala 201:45]
  assign _T_603 = legal_address & _T_515; // @[TLB.scala 197:19]
  assign prot_al = _T_603 | cacheable; // @[TLB.scala 202:46]
  assign _T_655 = $signed(_T_382) & 41'shca000000; // @[Parameters.scala 121:52]
  assign _T_656 = $signed(_T_655) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_667 = _T_656 | _T_553; // @[Parameters.scala 148:89]
  assign _T_668 = _T_667 | _T_558; // @[Parameters.scala 148:89]
  assign _T_675 = legal_address & _T_668; // @[TLB.scala 197:19]
  assign prot_x = _T_675 & pmp_io_x; // @[TLB.scala 204:40]
  assign _T_701 = $signed(_T_377) & 41'shca010000; // @[Parameters.scala 121:52]
  assign _T_702 = $signed(_T_701) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_706 = $signed(_T_382) & 41'shca012000; // @[Parameters.scala 121:52]
  assign _T_707 = $signed(_T_706) == 41'sh0; // @[Parameters.scala 121:67]
  assign _T_713 = _T_489 | _T_702; // @[Parameters.scala 148:89]
  assign _T_714 = _T_713 | _T_707; // @[Parameters.scala 148:89]
  assign _T_715 = _T_714 | _T_558; // @[Parameters.scala 148:89]
  assign prot_eff = legal_address & _T_715; // @[TLB.scala 197:19]
  assign _T_722 = sectored_entries_0_valid_0 | sectored_entries_0_valid_1; // @[package.scala 63:59]
  assign _T_723 = _T_722 | sectored_entries_0_valid_2; // @[package.scala 63:59]
  assign _T_724 = _T_723 | sectored_entries_0_valid_3; // @[package.scala 63:59]
  assign _T_725 = sectored_entries_0_tag ^ vpn; // @[TLB.scala 103:43]
  assign _T_727 = _T_725[26:2] == 25'h0; // @[TLB.scala 103:68]
  assign sector_hits_0 = _T_724 & _T_727; // @[TLB.scala 102:42]
  assign _T_728 = sectored_entries_1_valid_0 | sectored_entries_1_valid_1; // @[package.scala 63:59]
  assign _T_729 = _T_728 | sectored_entries_1_valid_2; // @[package.scala 63:59]
  assign _T_730 = _T_729 | sectored_entries_1_valid_3; // @[package.scala 63:59]
  assign _T_731 = sectored_entries_1_tag ^ vpn; // @[TLB.scala 103:43]
  assign _T_733 = _T_731[26:2] == 25'h0; // @[TLB.scala 103:68]
  assign sector_hits_1 = _T_730 & _T_733; // @[TLB.scala 102:42]
  assign _T_734 = sectored_entries_2_valid_0 | sectored_entries_2_valid_1; // @[package.scala 63:59]
  assign _T_735 = _T_734 | sectored_entries_2_valid_2; // @[package.scala 63:59]
  assign _T_736 = _T_735 | sectored_entries_2_valid_3; // @[package.scala 63:59]
  assign _T_737 = sectored_entries_2_tag ^ vpn; // @[TLB.scala 103:43]
  assign _T_739 = _T_737[26:2] == 25'h0; // @[TLB.scala 103:68]
  assign sector_hits_2 = _T_736 & _T_739; // @[TLB.scala 102:42]
  assign _T_740 = sectored_entries_3_valid_0 | sectored_entries_3_valid_1; // @[package.scala 63:59]
  assign _T_741 = _T_740 | sectored_entries_3_valid_2; // @[package.scala 63:59]
  assign _T_742 = _T_741 | sectored_entries_3_valid_3; // @[package.scala 63:59]
  assign _T_743 = sectored_entries_3_tag ^ vpn; // @[TLB.scala 103:43]
  assign _T_745 = _T_743[26:2] == 25'h0; // @[TLB.scala 103:68]
  assign sector_hits_3 = _T_742 & _T_745; // @[TLB.scala 102:42]
  assign _T_746 = sectored_entries_4_valid_0 | sectored_entries_4_valid_1; // @[package.scala 63:59]
  assign _T_747 = _T_746 | sectored_entries_4_valid_2; // @[package.scala 63:59]
  assign _T_748 = _T_747 | sectored_entries_4_valid_3; // @[package.scala 63:59]
  assign _T_749 = sectored_entries_4_tag ^ vpn; // @[TLB.scala 103:43]
  assign _T_751 = _T_749[26:2] == 25'h0; // @[TLB.scala 103:68]
  assign sector_hits_4 = _T_748 & _T_751; // @[TLB.scala 102:42]
  assign _T_752 = sectored_entries_5_valid_0 | sectored_entries_5_valid_1; // @[package.scala 63:59]
  assign _T_753 = _T_752 | sectored_entries_5_valid_2; // @[package.scala 63:59]
  assign _T_754 = _T_753 | sectored_entries_5_valid_3; // @[package.scala 63:59]
  assign _T_755 = sectored_entries_5_tag ^ vpn; // @[TLB.scala 103:43]
  assign _T_757 = _T_755[26:2] == 25'h0; // @[TLB.scala 103:68]
  assign sector_hits_5 = _T_754 & _T_757; // @[TLB.scala 102:42]
  assign _T_758 = sectored_entries_6_valid_0 | sectored_entries_6_valid_1; // @[package.scala 63:59]
  assign _T_759 = _T_758 | sectored_entries_6_valid_2; // @[package.scala 63:59]
  assign _T_760 = _T_759 | sectored_entries_6_valid_3; // @[package.scala 63:59]
  assign _T_761 = sectored_entries_6_tag ^ vpn; // @[TLB.scala 103:43]
  assign _T_763 = _T_761[26:2] == 25'h0; // @[TLB.scala 103:68]
  assign sector_hits_6 = _T_760 & _T_763; // @[TLB.scala 102:42]
  assign _T_764 = sectored_entries_7_valid_0 | sectored_entries_7_valid_1; // @[package.scala 63:59]
  assign _T_765 = _T_764 | sectored_entries_7_valid_2; // @[package.scala 63:59]
  assign _T_766 = _T_765 | sectored_entries_7_valid_3; // @[package.scala 63:59]
  assign _T_767 = sectored_entries_7_tag ^ vpn; // @[TLB.scala 103:43]
  assign _T_769 = _T_767[26:2] == 25'h0; // @[TLB.scala 103:68]
  assign sector_hits_7 = _T_766 & _T_769; // @[TLB.scala 102:42]
  assign _T_774 = superpage_entries_0_tag[26:18] == vpn[26:18]; // @[TLB.scala 110:79]
  assign _T_776 = superpage_entries_0_valid_0 & _T_774; // @[TLB.scala 110:31]
  assign _T_777 = superpage_entries_0_level < 2'h1; // @[TLB.scala 109:30]
  assign _T_781 = superpage_entries_0_tag[17:9] == vpn[17:9]; // @[TLB.scala 110:79]
  assign _T_782 = _T_777 | _T_781; // @[TLB.scala 110:42]
  assign superpage_hits_0 = _T_776 & _T_782; // @[TLB.scala 110:31]
  assign _T_794 = superpage_entries_1_tag[26:18] == vpn[26:18]; // @[TLB.scala 110:79]
  assign _T_796 = superpage_entries_1_valid_0 & _T_794; // @[TLB.scala 110:31]
  assign _T_797 = superpage_entries_1_level < 2'h1; // @[TLB.scala 109:30]
  assign _T_801 = superpage_entries_1_tag[17:9] == vpn[17:9]; // @[TLB.scala 110:79]
  assign _T_802 = _T_797 | _T_801; // @[TLB.scala 110:42]
  assign superpage_hits_1 = _T_796 & _T_802; // @[TLB.scala 110:31]
  assign _T_814 = superpage_entries_2_tag[26:18] == vpn[26:18]; // @[TLB.scala 110:79]
  assign _T_816 = superpage_entries_2_valid_0 & _T_814; // @[TLB.scala 110:31]
  assign _T_817 = superpage_entries_2_level < 2'h1; // @[TLB.scala 109:30]
  assign _T_821 = superpage_entries_2_tag[17:9] == vpn[17:9]; // @[TLB.scala 110:79]
  assign _T_822 = _T_817 | _T_821; // @[TLB.scala 110:42]
  assign superpage_hits_2 = _T_816 & _T_822; // @[TLB.scala 110:31]
  assign _T_834 = superpage_entries_3_tag[26:18] == vpn[26:18]; // @[TLB.scala 110:79]
  assign _T_836 = superpage_entries_3_valid_0 & _T_834; // @[TLB.scala 110:31]
  assign _T_837 = superpage_entries_3_level < 2'h1; // @[TLB.scala 109:30]
  assign _T_841 = superpage_entries_3_tag[17:9] == vpn[17:9]; // @[TLB.scala 110:79]
  assign _T_842 = _T_837 | _T_841; // @[TLB.scala 110:42]
  assign superpage_hits_3 = _T_836 & _T_842; // @[TLB.scala 110:31]
  assign _GEN_1 = 2'h1 == vpn[1:0] ? sectored_entries_0_valid_1 : sectored_entries_0_valid_0; // @[TLB.scala 115:20]
  assign _GEN_2 = 2'h2 == vpn[1:0] ? sectored_entries_0_valid_2 : _GEN_1; // @[TLB.scala 115:20]
  assign _GEN_3 = 2'h3 == vpn[1:0] ? sectored_entries_0_valid_3 : _GEN_2; // @[TLB.scala 115:20]
  assign _T_854 = _GEN_3 & _T_727; // @[TLB.scala 115:20]
  assign hitsVec_0 = vm_enabled & _T_854; // @[TLB.scala 209:44]
  assign _GEN_5 = 2'h1 == vpn[1:0] ? sectored_entries_1_valid_1 : sectored_entries_1_valid_0; // @[TLB.scala 115:20]
  assign _GEN_6 = 2'h2 == vpn[1:0] ? sectored_entries_1_valid_2 : _GEN_5; // @[TLB.scala 115:20]
  assign _GEN_7 = 2'h3 == vpn[1:0] ? sectored_entries_1_valid_3 : _GEN_6; // @[TLB.scala 115:20]
  assign _T_859 = _GEN_7 & _T_733; // @[TLB.scala 115:20]
  assign hitsVec_1 = vm_enabled & _T_859; // @[TLB.scala 209:44]
  assign _GEN_9 = 2'h1 == vpn[1:0] ? sectored_entries_2_valid_1 : sectored_entries_2_valid_0; // @[TLB.scala 115:20]
  assign _GEN_10 = 2'h2 == vpn[1:0] ? sectored_entries_2_valid_2 : _GEN_9; // @[TLB.scala 115:20]
  assign _GEN_11 = 2'h3 == vpn[1:0] ? sectored_entries_2_valid_3 : _GEN_10; // @[TLB.scala 115:20]
  assign _T_864 = _GEN_11 & _T_739; // @[TLB.scala 115:20]
  assign hitsVec_2 = vm_enabled & _T_864; // @[TLB.scala 209:44]
  assign _GEN_13 = 2'h1 == vpn[1:0] ? sectored_entries_3_valid_1 : sectored_entries_3_valid_0; // @[TLB.scala 115:20]
  assign _GEN_14 = 2'h2 == vpn[1:0] ? sectored_entries_3_valid_2 : _GEN_13; // @[TLB.scala 115:20]
  assign _GEN_15 = 2'h3 == vpn[1:0] ? sectored_entries_3_valid_3 : _GEN_14; // @[TLB.scala 115:20]
  assign _T_869 = _GEN_15 & _T_745; // @[TLB.scala 115:20]
  assign hitsVec_3 = vm_enabled & _T_869; // @[TLB.scala 209:44]
  assign _GEN_17 = 2'h1 == vpn[1:0] ? sectored_entries_4_valid_1 : sectored_entries_4_valid_0; // @[TLB.scala 115:20]
  assign _GEN_18 = 2'h2 == vpn[1:0] ? sectored_entries_4_valid_2 : _GEN_17; // @[TLB.scala 115:20]
  assign _GEN_19 = 2'h3 == vpn[1:0] ? sectored_entries_4_valid_3 : _GEN_18; // @[TLB.scala 115:20]
  assign _T_874 = _GEN_19 & _T_751; // @[TLB.scala 115:20]
  assign hitsVec_4 = vm_enabled & _T_874; // @[TLB.scala 209:44]
  assign _GEN_21 = 2'h1 == vpn[1:0] ? sectored_entries_5_valid_1 : sectored_entries_5_valid_0; // @[TLB.scala 115:20]
  assign _GEN_22 = 2'h2 == vpn[1:0] ? sectored_entries_5_valid_2 : _GEN_21; // @[TLB.scala 115:20]
  assign _GEN_23 = 2'h3 == vpn[1:0] ? sectored_entries_5_valid_3 : _GEN_22; // @[TLB.scala 115:20]
  assign _T_879 = _GEN_23 & _T_757; // @[TLB.scala 115:20]
  assign hitsVec_5 = vm_enabled & _T_879; // @[TLB.scala 209:44]
  assign _GEN_25 = 2'h1 == vpn[1:0] ? sectored_entries_6_valid_1 : sectored_entries_6_valid_0; // @[TLB.scala 115:20]
  assign _GEN_26 = 2'h2 == vpn[1:0] ? sectored_entries_6_valid_2 : _GEN_25; // @[TLB.scala 115:20]
  assign _GEN_27 = 2'h3 == vpn[1:0] ? sectored_entries_6_valid_3 : _GEN_26; // @[TLB.scala 115:20]
  assign _T_884 = _GEN_27 & _T_763; // @[TLB.scala 115:20]
  assign hitsVec_6 = vm_enabled & _T_884; // @[TLB.scala 209:44]
  assign _GEN_29 = 2'h1 == vpn[1:0] ? sectored_entries_7_valid_1 : sectored_entries_7_valid_0; // @[TLB.scala 115:20]
  assign _GEN_30 = 2'h2 == vpn[1:0] ? sectored_entries_7_valid_2 : _GEN_29; // @[TLB.scala 115:20]
  assign _GEN_31 = 2'h3 == vpn[1:0] ? sectored_entries_7_valid_3 : _GEN_30; // @[TLB.scala 115:20]
  assign _T_889 = _GEN_31 & _T_769; // @[TLB.scala 115:20]
  assign hitsVec_7 = vm_enabled & _T_889; // @[TLB.scala 209:44]
  assign hitsVec_8 = vm_enabled & superpage_hits_0; // @[TLB.scala 209:44]
  assign hitsVec_9 = vm_enabled & superpage_hits_1; // @[TLB.scala 209:44]
  assign hitsVec_10 = vm_enabled & superpage_hits_2; // @[TLB.scala 209:44]
  assign hitsVec_11 = vm_enabled & superpage_hits_3; // @[TLB.scala 209:44]
  assign _T_978 = special_entry_tag[26:18] == vpn[26:18]; // @[TLB.scala 110:79]
  assign _T_980 = special_entry_valid_0 & _T_978; // @[TLB.scala 110:31]
  assign _T_985 = special_entry_tag[17:9] == vpn[17:9]; // @[TLB.scala 110:79]
  assign _T_986 = _T_348 | _T_985; // @[TLB.scala 110:42]
  assign _T_987 = _T_980 & _T_986; // @[TLB.scala 110:31]
  assign _T_992 = special_entry_tag[8:0] == vpn[8:0]; // @[TLB.scala 110:79]
  assign _T_993 = _T_354 | _T_992; // @[TLB.scala 110:42]
  assign _T_994 = _T_987 & _T_993; // @[TLB.scala 110:31]
  assign hitsVec_12 = vm_enabled & _T_994; // @[TLB.scala 209:44]
  assign _T_999 = {hitsVec_5,hitsVec_4,hitsVec_3,hitsVec_2,hitsVec_1,hitsVec_0}; // @[Cat.scala 30:58]
  assign real_hits = {hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,_T_999}; // @[Cat.scala 30:58]
  assign hits = {~vm_enabled,hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,_T_999}; // @[Cat.scala 30:58]
  assign _GEN_33 = 2'h1 == vpn[1:0] ? sectored_entries_0_data_1 : sectored_entries_0_data_0;
  assign _GEN_34 = 2'h2 == vpn[1:0] ? sectored_entries_0_data_2 : _GEN_33;
  assign _GEN_35 = 2'h3 == vpn[1:0] ? sectored_entries_0_data_3 : _GEN_34;
  assign _GEN_37 = 2'h1 == vpn[1:0] ? sectored_entries_1_data_1 : sectored_entries_1_data_0;
  assign _GEN_38 = 2'h2 == vpn[1:0] ? sectored_entries_1_data_2 : _GEN_37;
  assign _GEN_39 = 2'h3 == vpn[1:0] ? sectored_entries_1_data_3 : _GEN_38;
  assign _GEN_41 = 2'h1 == vpn[1:0] ? sectored_entries_2_data_1 : sectored_entries_2_data_0;
  assign _GEN_42 = 2'h2 == vpn[1:0] ? sectored_entries_2_data_2 : _GEN_41;
  assign _GEN_43 = 2'h3 == vpn[1:0] ? sectored_entries_2_data_3 : _GEN_42;
  assign _GEN_45 = 2'h1 == vpn[1:0] ? sectored_entries_3_data_1 : sectored_entries_3_data_0;
  assign _GEN_46 = 2'h2 == vpn[1:0] ? sectored_entries_3_data_2 : _GEN_45;
  assign _GEN_47 = 2'h3 == vpn[1:0] ? sectored_entries_3_data_3 : _GEN_46;
  assign _GEN_49 = 2'h1 == vpn[1:0] ? sectored_entries_4_data_1 : sectored_entries_4_data_0;
  assign _GEN_50 = 2'h2 == vpn[1:0] ? sectored_entries_4_data_2 : _GEN_49;
  assign _GEN_51 = 2'h3 == vpn[1:0] ? sectored_entries_4_data_3 : _GEN_50;
  assign _GEN_53 = 2'h1 == vpn[1:0] ? sectored_entries_5_data_1 : sectored_entries_5_data_0;
  assign _GEN_54 = 2'h2 == vpn[1:0] ? sectored_entries_5_data_2 : _GEN_53;
  assign _GEN_55 = 2'h3 == vpn[1:0] ? sectored_entries_5_data_3 : _GEN_54;
  assign _GEN_57 = 2'h1 == vpn[1:0] ? sectored_entries_6_data_1 : sectored_entries_6_data_0;
  assign _GEN_58 = 2'h2 == vpn[1:0] ? sectored_entries_6_data_2 : _GEN_57;
  assign _GEN_59 = 2'h3 == vpn[1:0] ? sectored_entries_6_data_3 : _GEN_58;
  assign _GEN_61 = 2'h1 == vpn[1:0] ? sectored_entries_7_data_1 : sectored_entries_7_data_0;
  assign _GEN_62 = 2'h2 == vpn[1:0] ? sectored_entries_7_data_2 : _GEN_61;
  assign _GEN_63 = 2'h3 == vpn[1:0] ? sectored_entries_7_data_3 : _GEN_62;
  assign _T_1199 = _T_777 ? vpn : 27'h0; // @[TLB.scala 124:30]
  assign _GEN_956 = {{7'd0}, superpage_entries_0_data_0[33:14]}; // @[TLB.scala 124:49]
  assign _T_1200 = _T_1199 | _GEN_956; // @[TLB.scala 124:49]
  assign _T_1206 = vpn | _GEN_956; // @[TLB.scala 124:49]
  assign _T_1208 = {superpage_entries_0_data_0[33:32],_T_1200[17:9],_T_1206[8:0]}; // @[Cat.scala 30:58]
  assign _T_1232 = _T_797 ? vpn : 27'h0; // @[TLB.scala 124:30]
  assign _GEN_958 = {{7'd0}, superpage_entries_1_data_0[33:14]}; // @[TLB.scala 124:49]
  assign _T_1233 = _T_1232 | _GEN_958; // @[TLB.scala 124:49]
  assign _T_1239 = vpn | _GEN_958; // @[TLB.scala 124:49]
  assign _T_1241 = {superpage_entries_1_data_0[33:32],_T_1233[17:9],_T_1239[8:0]}; // @[Cat.scala 30:58]
  assign _T_1265 = _T_817 ? vpn : 27'h0; // @[TLB.scala 124:30]
  assign _GEN_960 = {{7'd0}, superpage_entries_2_data_0[33:14]}; // @[TLB.scala 124:49]
  assign _T_1266 = _T_1265 | _GEN_960; // @[TLB.scala 124:49]
  assign _T_1272 = vpn | _GEN_960; // @[TLB.scala 124:49]
  assign _T_1274 = {superpage_entries_2_data_0[33:32],_T_1266[17:9],_T_1272[8:0]}; // @[Cat.scala 30:58]
  assign _T_1298 = _T_837 ? vpn : 27'h0; // @[TLB.scala 124:30]
  assign _GEN_962 = {{7'd0}, superpage_entries_3_data_0[33:14]}; // @[TLB.scala 124:49]
  assign _T_1299 = _T_1298 | _GEN_962; // @[TLB.scala 124:49]
  assign _T_1305 = vpn | _GEN_962; // @[TLB.scala 124:49]
  assign _T_1307 = {superpage_entries_3_data_0[33:32],_T_1299[17:9],_T_1305[8:0]}; // @[Cat.scala 30:58]
  assign _T_1343 = hitsVec_0 ? _GEN_35[33:14] : 20'h0; // @[Mux.scala 19:72]
  assign _T_1344 = hitsVec_1 ? _GEN_39[33:14] : 20'h0; // @[Mux.scala 19:72]
  assign _T_1345 = hitsVec_2 ? _GEN_43[33:14] : 20'h0; // @[Mux.scala 19:72]
  assign _T_1346 = hitsVec_3 ? _GEN_47[33:14] : 20'h0; // @[Mux.scala 19:72]
  assign _T_1347 = hitsVec_4 ? _GEN_51[33:14] : 20'h0; // @[Mux.scala 19:72]
  assign _T_1348 = hitsVec_5 ? _GEN_55[33:14] : 20'h0; // @[Mux.scala 19:72]
  assign _T_1349 = hitsVec_6 ? _GEN_59[33:14] : 20'h0; // @[Mux.scala 19:72]
  assign _T_1350 = hitsVec_7 ? _GEN_63[33:14] : 20'h0; // @[Mux.scala 19:72]
  assign _T_1351 = hitsVec_8 ? _T_1208 : 20'h0; // @[Mux.scala 19:72]
  assign _T_1352 = hitsVec_9 ? _T_1241 : 20'h0; // @[Mux.scala 19:72]
  assign _T_1353 = hitsVec_10 ? _T_1274 : 20'h0; // @[Mux.scala 19:72]
  assign _T_1354 = hitsVec_11 ? _T_1307 : 20'h0; // @[Mux.scala 19:72]
  assign _T_1355 = hitsVec_12 ? _T_359 : 20'h0; // @[Mux.scala 19:72]
  assign _T_1356 = vm_enabled ? 20'h0 : vpn[19:0]; // @[Mux.scala 19:72]
  assign _T_1357 = _T_1343 | _T_1344; // @[Mux.scala 19:72]
  assign _T_1358 = _T_1357 | _T_1345; // @[Mux.scala 19:72]
  assign _T_1359 = _T_1358 | _T_1346; // @[Mux.scala 19:72]
  assign _T_1360 = _T_1359 | _T_1347; // @[Mux.scala 19:72]
  assign _T_1361 = _T_1360 | _T_1348; // @[Mux.scala 19:72]
  assign _T_1362 = _T_1361 | _T_1349; // @[Mux.scala 19:72]
  assign _T_1363 = _T_1362 | _T_1350; // @[Mux.scala 19:72]
  assign _T_1364 = _T_1363 | _T_1351; // @[Mux.scala 19:72]
  assign _T_1365 = _T_1364 | _T_1352; // @[Mux.scala 19:72]
  assign _T_1366 = _T_1365 | _T_1353; // @[Mux.scala 19:72]
  assign _T_1367 = _T_1366 | _T_1354; // @[Mux.scala 19:72]
  assign _T_1368 = _T_1367 | _T_1355; // @[Mux.scala 19:72]
  assign ppn = _T_1368 | _T_1356; // @[Mux.scala 19:72]
  assign _T_1385 = io_ptw_resp_valid & ~invalidate_refill; // @[TLB.scala 224:17]
  assign _GEN_966 = {{27'd0}, vpoffset_cfg_value}; // @[TLB.scala 227:31]
  assign _T_1387 = io_ptw_resp_bits_pte_ppn + _GEN_966; // @[TLB.scala 227:31]
  assign _T_1391 = io_ptw_resp_bits_pte_x & ~io_ptw_resp_bits_pte_w; // @[PTW.scala 77:44]
  assign _T_1392 = io_ptw_resp_bits_pte_r | _T_1391; // @[PTW.scala 77:38]
  assign _T_1393 = io_ptw_resp_bits_pte_v & _T_1392; // @[PTW.scala 77:32]
  assign _T_1394 = _T_1393 & io_ptw_resp_bits_pte_a; // @[PTW.scala 77:52]
  assign _T_1395 = _T_1394 & io_ptw_resp_bits_pte_r; // @[PTW.scala 81:35]
  assign _T_1401 = _T_1394 & io_ptw_resp_bits_pte_w; // @[PTW.scala 82:35]
  assign _T_1402 = _T_1401 & io_ptw_resp_bits_pte_d; // @[PTW.scala 82:40]
  assign _T_1403 = vpoffset_cfg_value == 27'h0; // @[TLB.scala 231:55]
  assign _T_1404 = io_ptw_resp_bits_pte_u | _T_1403; // @[TLB.scala 231:32]
  assign _T_1405 = io_ptw_resp_bits_level != 2'h2; // @[TLB.scala 231:90]
  assign _T_1406 = _T_1404 | _T_1405; // @[TLB.scala 231:64]
  assign _T_1412 = _T_1394 & io_ptw_resp_bits_pte_x; // @[PTW.scala 83:35]
  assign _GEN_967 = {{27'd0}, requestedVPN}; // @[TLB.scala 231:133]
  assign _T_1413 = _T_1387 == _GEN_967; // @[TLB.scala 231:133]
  assign _T_1420 = _T_1413 & _T_1412; // @[TLB.scala 231:120]
  assign _T_1421 = _T_1406 ? _T_1412 : _T_1420; // @[TLB.scala 231:25]
  assign _T_1430 = {prot_x,prot_r,prot_al,prot_al,prot_eff,cacheable,1'h0}; // @[TLB.scala 138:26]
  assign _T_1438 = {refill_ppn,io_ptw_resp_bits_pte_u,io_ptw_resp_bits_pte_g,io_ptw_resp_bits_ae,_T_1402,_T_1421,_T_1395,prot_w,_T_1430}; // @[TLB.scala 138:26]
  assign _T_1439 = io_ptw_resp_bits_level < 2'h2; // @[TLB.scala 253:40]
  assign _T_1440 = r_superpage_repl_addr == 2'h0; // @[TLB.scala 254:82]
  assign _GEN_67 = _T_1440 | superpage_entries_0_valid_0; // @[TLB.scala 254:89]
  assign _T_1456 = r_superpage_repl_addr == 2'h1; // @[TLB.scala 254:82]
  assign _GEN_71 = _T_1456 | superpage_entries_1_valid_0; // @[TLB.scala 254:89]
  assign _T_1472 = r_superpage_repl_addr == 2'h2; // @[TLB.scala 254:82]
  assign _GEN_75 = _T_1472 | superpage_entries_2_valid_0; // @[TLB.scala 254:89]
  assign _T_1488 = r_superpage_repl_addr == 2'h3; // @[TLB.scala 254:82]
  assign _GEN_79 = _T_1488 | superpage_entries_3_valid_0; // @[TLB.scala 254:89]
  assign _T_1504 = r_sectored_hit ? r_sectored_hit_addr : r_sectored_repl_addr; // @[TLB.scala 258:22]
  assign _T_1505 = _T_1504 == 3'h0; // @[TLB.scala 259:65]
  assign _GEN_81 = r_sectored_hit ? sectored_entries_0_valid_0 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_82 = r_sectored_hit ? sectored_entries_0_valid_1 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_83 = r_sectored_hit ? sectored_entries_0_valid_2 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_84 = r_sectored_hit ? sectored_entries_0_valid_3 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_968 = 2'h0 == r_refill_tag[1:0]; // @[TLB.scala 137:18]
  assign _GEN_85 = _GEN_968 | _GEN_81; // @[TLB.scala 137:18]
  assign _GEN_969 = 2'h1 == r_refill_tag[1:0]; // @[TLB.scala 137:18]
  assign _GEN_86 = _GEN_969 | _GEN_82; // @[TLB.scala 137:18]
  assign _GEN_970 = 2'h2 == r_refill_tag[1:0]; // @[TLB.scala 137:18]
  assign _GEN_87 = _GEN_970 | _GEN_83; // @[TLB.scala 137:18]
  assign _GEN_971 = 2'h3 == r_refill_tag[1:0]; // @[TLB.scala 137:18]
  assign _GEN_88 = _GEN_971 | _GEN_84; // @[TLB.scala 137:18]
  assign _GEN_93 = _T_1505 ? _GEN_85 : sectored_entries_0_valid_0; // @[TLB.scala 259:72]
  assign _GEN_94 = _T_1505 ? _GEN_86 : sectored_entries_0_valid_1; // @[TLB.scala 259:72]
  assign _GEN_95 = _T_1505 ? _GEN_87 : sectored_entries_0_valid_2; // @[TLB.scala 259:72]
  assign _GEN_96 = _T_1505 ? _GEN_88 : sectored_entries_0_valid_3; // @[TLB.scala 259:72]
  assign _T_1522 = _T_1504 == 3'h1; // @[TLB.scala 259:65]
  assign _GEN_103 = r_sectored_hit ? sectored_entries_1_valid_0 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_104 = r_sectored_hit ? sectored_entries_1_valid_1 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_105 = r_sectored_hit ? sectored_entries_1_valid_2 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_106 = r_sectored_hit ? sectored_entries_1_valid_3 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_107 = _GEN_968 | _GEN_103; // @[TLB.scala 137:18]
  assign _GEN_108 = _GEN_969 | _GEN_104; // @[TLB.scala 137:18]
  assign _GEN_109 = _GEN_970 | _GEN_105; // @[TLB.scala 137:18]
  assign _GEN_110 = _GEN_971 | _GEN_106; // @[TLB.scala 137:18]
  assign _GEN_115 = _T_1522 ? _GEN_107 : sectored_entries_1_valid_0; // @[TLB.scala 259:72]
  assign _GEN_116 = _T_1522 ? _GEN_108 : sectored_entries_1_valid_1; // @[TLB.scala 259:72]
  assign _GEN_117 = _T_1522 ? _GEN_109 : sectored_entries_1_valid_2; // @[TLB.scala 259:72]
  assign _GEN_118 = _T_1522 ? _GEN_110 : sectored_entries_1_valid_3; // @[TLB.scala 259:72]
  assign _T_1539 = _T_1504 == 3'h2; // @[TLB.scala 259:65]
  assign _GEN_125 = r_sectored_hit ? sectored_entries_2_valid_0 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_126 = r_sectored_hit ? sectored_entries_2_valid_1 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_127 = r_sectored_hit ? sectored_entries_2_valid_2 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_128 = r_sectored_hit ? sectored_entries_2_valid_3 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_129 = _GEN_968 | _GEN_125; // @[TLB.scala 137:18]
  assign _GEN_130 = _GEN_969 | _GEN_126; // @[TLB.scala 137:18]
  assign _GEN_131 = _GEN_970 | _GEN_127; // @[TLB.scala 137:18]
  assign _GEN_132 = _GEN_971 | _GEN_128; // @[TLB.scala 137:18]
  assign _GEN_137 = _T_1539 ? _GEN_129 : sectored_entries_2_valid_0; // @[TLB.scala 259:72]
  assign _GEN_138 = _T_1539 ? _GEN_130 : sectored_entries_2_valid_1; // @[TLB.scala 259:72]
  assign _GEN_139 = _T_1539 ? _GEN_131 : sectored_entries_2_valid_2; // @[TLB.scala 259:72]
  assign _GEN_140 = _T_1539 ? _GEN_132 : sectored_entries_2_valid_3; // @[TLB.scala 259:72]
  assign _T_1556 = _T_1504 == 3'h3; // @[TLB.scala 259:65]
  assign _GEN_147 = r_sectored_hit ? sectored_entries_3_valid_0 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_148 = r_sectored_hit ? sectored_entries_3_valid_1 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_149 = r_sectored_hit ? sectored_entries_3_valid_2 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_150 = r_sectored_hit ? sectored_entries_3_valid_3 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_151 = _GEN_968 | _GEN_147; // @[TLB.scala 137:18]
  assign _GEN_152 = _GEN_969 | _GEN_148; // @[TLB.scala 137:18]
  assign _GEN_153 = _GEN_970 | _GEN_149; // @[TLB.scala 137:18]
  assign _GEN_154 = _GEN_971 | _GEN_150; // @[TLB.scala 137:18]
  assign _GEN_159 = _T_1556 ? _GEN_151 : sectored_entries_3_valid_0; // @[TLB.scala 259:72]
  assign _GEN_160 = _T_1556 ? _GEN_152 : sectored_entries_3_valid_1; // @[TLB.scala 259:72]
  assign _GEN_161 = _T_1556 ? _GEN_153 : sectored_entries_3_valid_2; // @[TLB.scala 259:72]
  assign _GEN_162 = _T_1556 ? _GEN_154 : sectored_entries_3_valid_3; // @[TLB.scala 259:72]
  assign _T_1573 = _T_1504 == 3'h4; // @[TLB.scala 259:65]
  assign _GEN_169 = r_sectored_hit ? sectored_entries_4_valid_0 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_170 = r_sectored_hit ? sectored_entries_4_valid_1 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_171 = r_sectored_hit ? sectored_entries_4_valid_2 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_172 = r_sectored_hit ? sectored_entries_4_valid_3 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_173 = _GEN_968 | _GEN_169; // @[TLB.scala 137:18]
  assign _GEN_174 = _GEN_969 | _GEN_170; // @[TLB.scala 137:18]
  assign _GEN_175 = _GEN_970 | _GEN_171; // @[TLB.scala 137:18]
  assign _GEN_176 = _GEN_971 | _GEN_172; // @[TLB.scala 137:18]
  assign _GEN_181 = _T_1573 ? _GEN_173 : sectored_entries_4_valid_0; // @[TLB.scala 259:72]
  assign _GEN_182 = _T_1573 ? _GEN_174 : sectored_entries_4_valid_1; // @[TLB.scala 259:72]
  assign _GEN_183 = _T_1573 ? _GEN_175 : sectored_entries_4_valid_2; // @[TLB.scala 259:72]
  assign _GEN_184 = _T_1573 ? _GEN_176 : sectored_entries_4_valid_3; // @[TLB.scala 259:72]
  assign _T_1590 = _T_1504 == 3'h5; // @[TLB.scala 259:65]
  assign _GEN_191 = r_sectored_hit ? sectored_entries_5_valid_0 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_192 = r_sectored_hit ? sectored_entries_5_valid_1 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_193 = r_sectored_hit ? sectored_entries_5_valid_2 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_194 = r_sectored_hit ? sectored_entries_5_valid_3 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_195 = _GEN_968 | _GEN_191; // @[TLB.scala 137:18]
  assign _GEN_196 = _GEN_969 | _GEN_192; // @[TLB.scala 137:18]
  assign _GEN_197 = _GEN_970 | _GEN_193; // @[TLB.scala 137:18]
  assign _GEN_198 = _GEN_971 | _GEN_194; // @[TLB.scala 137:18]
  assign _GEN_203 = _T_1590 ? _GEN_195 : sectored_entries_5_valid_0; // @[TLB.scala 259:72]
  assign _GEN_204 = _T_1590 ? _GEN_196 : sectored_entries_5_valid_1; // @[TLB.scala 259:72]
  assign _GEN_205 = _T_1590 ? _GEN_197 : sectored_entries_5_valid_2; // @[TLB.scala 259:72]
  assign _GEN_206 = _T_1590 ? _GEN_198 : sectored_entries_5_valid_3; // @[TLB.scala 259:72]
  assign _T_1607 = _T_1504 == 3'h6; // @[TLB.scala 259:65]
  assign _GEN_213 = r_sectored_hit ? sectored_entries_6_valid_0 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_214 = r_sectored_hit ? sectored_entries_6_valid_1 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_215 = r_sectored_hit ? sectored_entries_6_valid_2 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_216 = r_sectored_hit ? sectored_entries_6_valid_3 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_217 = _GEN_968 | _GEN_213; // @[TLB.scala 137:18]
  assign _GEN_218 = _GEN_969 | _GEN_214; // @[TLB.scala 137:18]
  assign _GEN_219 = _GEN_970 | _GEN_215; // @[TLB.scala 137:18]
  assign _GEN_220 = _GEN_971 | _GEN_216; // @[TLB.scala 137:18]
  assign _GEN_225 = _T_1607 ? _GEN_217 : sectored_entries_6_valid_0; // @[TLB.scala 259:72]
  assign _GEN_226 = _T_1607 ? _GEN_218 : sectored_entries_6_valid_1; // @[TLB.scala 259:72]
  assign _GEN_227 = _T_1607 ? _GEN_219 : sectored_entries_6_valid_2; // @[TLB.scala 259:72]
  assign _GEN_228 = _T_1607 ? _GEN_220 : sectored_entries_6_valid_3; // @[TLB.scala 259:72]
  assign _T_1624 = _T_1504 == 3'h7; // @[TLB.scala 259:65]
  assign _GEN_235 = r_sectored_hit ? sectored_entries_7_valid_0 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_236 = r_sectored_hit ? sectored_entries_7_valid_1 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_237 = r_sectored_hit ? sectored_entries_7_valid_2 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_238 = r_sectored_hit ? sectored_entries_7_valid_3 : 1'h0; // @[TLB.scala 260:32]
  assign _GEN_239 = _GEN_968 | _GEN_235; // @[TLB.scala 137:18]
  assign _GEN_240 = _GEN_969 | _GEN_236; // @[TLB.scala 137:18]
  assign _GEN_241 = _GEN_970 | _GEN_237; // @[TLB.scala 137:18]
  assign _GEN_242 = _GEN_971 | _GEN_238; // @[TLB.scala 137:18]
  assign _GEN_247 = _T_1624 ? _GEN_239 : sectored_entries_7_valid_0; // @[TLB.scala 259:72]
  assign _GEN_248 = _T_1624 ? _GEN_240 : sectored_entries_7_valid_1; // @[TLB.scala 259:72]
  assign _GEN_249 = _T_1624 ? _GEN_241 : sectored_entries_7_valid_2; // @[TLB.scala 259:72]
  assign _GEN_250 = _T_1624 ? _GEN_242 : sectored_entries_7_valid_3; // @[TLB.scala 259:72]
  assign _GEN_259 = _T_1439 ? _GEN_67 : superpage_entries_0_valid_0; // @[TLB.scala 253:54]
  assign _GEN_263 = _T_1439 ? _GEN_71 : superpage_entries_1_valid_0; // @[TLB.scala 253:54]
  assign _GEN_267 = _T_1439 ? _GEN_75 : superpage_entries_2_valid_0; // @[TLB.scala 253:54]
  assign _GEN_271 = _T_1439 ? _GEN_79 : superpage_entries_3_valid_0; // @[TLB.scala 253:54]
  assign _GEN_273 = _T_1439 ? sectored_entries_0_valid_0 : _GEN_93; // @[TLB.scala 253:54]
  assign _GEN_274 = _T_1439 ? sectored_entries_0_valid_1 : _GEN_94; // @[TLB.scala 253:54]
  assign _GEN_275 = _T_1439 ? sectored_entries_0_valid_2 : _GEN_95; // @[TLB.scala 253:54]
  assign _GEN_276 = _T_1439 ? sectored_entries_0_valid_3 : _GEN_96; // @[TLB.scala 253:54]
  assign _GEN_283 = _T_1439 ? sectored_entries_1_valid_0 : _GEN_115; // @[TLB.scala 253:54]
  assign _GEN_284 = _T_1439 ? sectored_entries_1_valid_1 : _GEN_116; // @[TLB.scala 253:54]
  assign _GEN_285 = _T_1439 ? sectored_entries_1_valid_2 : _GEN_117; // @[TLB.scala 253:54]
  assign _GEN_286 = _T_1439 ? sectored_entries_1_valid_3 : _GEN_118; // @[TLB.scala 253:54]
  assign _GEN_293 = _T_1439 ? sectored_entries_2_valid_0 : _GEN_137; // @[TLB.scala 253:54]
  assign _GEN_294 = _T_1439 ? sectored_entries_2_valid_1 : _GEN_138; // @[TLB.scala 253:54]
  assign _GEN_295 = _T_1439 ? sectored_entries_2_valid_2 : _GEN_139; // @[TLB.scala 253:54]
  assign _GEN_296 = _T_1439 ? sectored_entries_2_valid_3 : _GEN_140; // @[TLB.scala 253:54]
  assign _GEN_303 = _T_1439 ? sectored_entries_3_valid_0 : _GEN_159; // @[TLB.scala 253:54]
  assign _GEN_304 = _T_1439 ? sectored_entries_3_valid_1 : _GEN_160; // @[TLB.scala 253:54]
  assign _GEN_305 = _T_1439 ? sectored_entries_3_valid_2 : _GEN_161; // @[TLB.scala 253:54]
  assign _GEN_306 = _T_1439 ? sectored_entries_3_valid_3 : _GEN_162; // @[TLB.scala 253:54]
  assign _GEN_313 = _T_1439 ? sectored_entries_4_valid_0 : _GEN_181; // @[TLB.scala 253:54]
  assign _GEN_314 = _T_1439 ? sectored_entries_4_valid_1 : _GEN_182; // @[TLB.scala 253:54]
  assign _GEN_315 = _T_1439 ? sectored_entries_4_valid_2 : _GEN_183; // @[TLB.scala 253:54]
  assign _GEN_316 = _T_1439 ? sectored_entries_4_valid_3 : _GEN_184; // @[TLB.scala 253:54]
  assign _GEN_323 = _T_1439 ? sectored_entries_5_valid_0 : _GEN_203; // @[TLB.scala 253:54]
  assign _GEN_324 = _T_1439 ? sectored_entries_5_valid_1 : _GEN_204; // @[TLB.scala 253:54]
  assign _GEN_325 = _T_1439 ? sectored_entries_5_valid_2 : _GEN_205; // @[TLB.scala 253:54]
  assign _GEN_326 = _T_1439 ? sectored_entries_5_valid_3 : _GEN_206; // @[TLB.scala 253:54]
  assign _GEN_333 = _T_1439 ? sectored_entries_6_valid_0 : _GEN_225; // @[TLB.scala 253:54]
  assign _GEN_334 = _T_1439 ? sectored_entries_6_valid_1 : _GEN_226; // @[TLB.scala 253:54]
  assign _GEN_335 = _T_1439 ? sectored_entries_6_valid_2 : _GEN_227; // @[TLB.scala 253:54]
  assign _GEN_336 = _T_1439 ? sectored_entries_6_valid_3 : _GEN_228; // @[TLB.scala 253:54]
  assign _GEN_343 = _T_1439 ? sectored_entries_7_valid_0 : _GEN_247; // @[TLB.scala 253:54]
  assign _GEN_344 = _T_1439 ? sectored_entries_7_valid_1 : _GEN_248; // @[TLB.scala 253:54]
  assign _GEN_345 = _T_1439 ? sectored_entries_7_valid_2 : _GEN_249; // @[TLB.scala 253:54]
  assign _GEN_346 = _T_1439 ? sectored_entries_7_valid_3 : _GEN_250; // @[TLB.scala 253:54]
  assign _GEN_355 = ~io_ptw_resp_bits_homogeneous | special_entry_valid_0; // @[TLB.scala 251:68]
  assign _GEN_359 = io_ptw_resp_bits_homogeneous ? _GEN_259 : superpage_entries_0_valid_0; // @[TLB.scala 251:68]
  assign _GEN_363 = io_ptw_resp_bits_homogeneous ? _GEN_263 : superpage_entries_1_valid_0; // @[TLB.scala 251:68]
  assign _GEN_367 = io_ptw_resp_bits_homogeneous ? _GEN_267 : superpage_entries_2_valid_0; // @[TLB.scala 251:68]
  assign _GEN_371 = io_ptw_resp_bits_homogeneous ? _GEN_271 : superpage_entries_3_valid_0; // @[TLB.scala 251:68]
  assign _GEN_373 = io_ptw_resp_bits_homogeneous ? _GEN_273 : sectored_entries_0_valid_0; // @[TLB.scala 251:68]
  assign _GEN_374 = io_ptw_resp_bits_homogeneous ? _GEN_274 : sectored_entries_0_valid_1; // @[TLB.scala 251:68]
  assign _GEN_375 = io_ptw_resp_bits_homogeneous ? _GEN_275 : sectored_entries_0_valid_2; // @[TLB.scala 251:68]
  assign _GEN_376 = io_ptw_resp_bits_homogeneous ? _GEN_276 : sectored_entries_0_valid_3; // @[TLB.scala 251:68]
  assign _GEN_383 = io_ptw_resp_bits_homogeneous ? _GEN_283 : sectored_entries_1_valid_0; // @[TLB.scala 251:68]
  assign _GEN_384 = io_ptw_resp_bits_homogeneous ? _GEN_284 : sectored_entries_1_valid_1; // @[TLB.scala 251:68]
  assign _GEN_385 = io_ptw_resp_bits_homogeneous ? _GEN_285 : sectored_entries_1_valid_2; // @[TLB.scala 251:68]
  assign _GEN_386 = io_ptw_resp_bits_homogeneous ? _GEN_286 : sectored_entries_1_valid_3; // @[TLB.scala 251:68]
  assign _GEN_393 = io_ptw_resp_bits_homogeneous ? _GEN_293 : sectored_entries_2_valid_0; // @[TLB.scala 251:68]
  assign _GEN_394 = io_ptw_resp_bits_homogeneous ? _GEN_294 : sectored_entries_2_valid_1; // @[TLB.scala 251:68]
  assign _GEN_395 = io_ptw_resp_bits_homogeneous ? _GEN_295 : sectored_entries_2_valid_2; // @[TLB.scala 251:68]
  assign _GEN_396 = io_ptw_resp_bits_homogeneous ? _GEN_296 : sectored_entries_2_valid_3; // @[TLB.scala 251:68]
  assign _GEN_403 = io_ptw_resp_bits_homogeneous ? _GEN_303 : sectored_entries_3_valid_0; // @[TLB.scala 251:68]
  assign _GEN_404 = io_ptw_resp_bits_homogeneous ? _GEN_304 : sectored_entries_3_valid_1; // @[TLB.scala 251:68]
  assign _GEN_405 = io_ptw_resp_bits_homogeneous ? _GEN_305 : sectored_entries_3_valid_2; // @[TLB.scala 251:68]
  assign _GEN_406 = io_ptw_resp_bits_homogeneous ? _GEN_306 : sectored_entries_3_valid_3; // @[TLB.scala 251:68]
  assign _GEN_413 = io_ptw_resp_bits_homogeneous ? _GEN_313 : sectored_entries_4_valid_0; // @[TLB.scala 251:68]
  assign _GEN_414 = io_ptw_resp_bits_homogeneous ? _GEN_314 : sectored_entries_4_valid_1; // @[TLB.scala 251:68]
  assign _GEN_415 = io_ptw_resp_bits_homogeneous ? _GEN_315 : sectored_entries_4_valid_2; // @[TLB.scala 251:68]
  assign _GEN_416 = io_ptw_resp_bits_homogeneous ? _GEN_316 : sectored_entries_4_valid_3; // @[TLB.scala 251:68]
  assign _GEN_423 = io_ptw_resp_bits_homogeneous ? _GEN_323 : sectored_entries_5_valid_0; // @[TLB.scala 251:68]
  assign _GEN_424 = io_ptw_resp_bits_homogeneous ? _GEN_324 : sectored_entries_5_valid_1; // @[TLB.scala 251:68]
  assign _GEN_425 = io_ptw_resp_bits_homogeneous ? _GEN_325 : sectored_entries_5_valid_2; // @[TLB.scala 251:68]
  assign _GEN_426 = io_ptw_resp_bits_homogeneous ? _GEN_326 : sectored_entries_5_valid_3; // @[TLB.scala 251:68]
  assign _GEN_433 = io_ptw_resp_bits_homogeneous ? _GEN_333 : sectored_entries_6_valid_0; // @[TLB.scala 251:68]
  assign _GEN_434 = io_ptw_resp_bits_homogeneous ? _GEN_334 : sectored_entries_6_valid_1; // @[TLB.scala 251:68]
  assign _GEN_435 = io_ptw_resp_bits_homogeneous ? _GEN_335 : sectored_entries_6_valid_2; // @[TLB.scala 251:68]
  assign _GEN_436 = io_ptw_resp_bits_homogeneous ? _GEN_336 : sectored_entries_6_valid_3; // @[TLB.scala 251:68]
  assign _GEN_443 = io_ptw_resp_bits_homogeneous ? _GEN_343 : sectored_entries_7_valid_0; // @[TLB.scala 251:68]
  assign _GEN_444 = io_ptw_resp_bits_homogeneous ? _GEN_344 : sectored_entries_7_valid_1; // @[TLB.scala 251:68]
  assign _GEN_445 = io_ptw_resp_bits_homogeneous ? _GEN_345 : sectored_entries_7_valid_2; // @[TLB.scala 251:68]
  assign _GEN_446 = io_ptw_resp_bits_homogeneous ? _GEN_346 : sectored_entries_7_valid_3; // @[TLB.scala 251:68]
  assign _GEN_455 = _T_1385 ? _GEN_355 : special_entry_valid_0; // @[TLB.scala 224:40]
  assign _GEN_459 = _T_1385 ? _GEN_359 : superpage_entries_0_valid_0; // @[TLB.scala 224:40]
  assign _GEN_463 = _T_1385 ? _GEN_363 : superpage_entries_1_valid_0; // @[TLB.scala 224:40]
  assign _GEN_467 = _T_1385 ? _GEN_367 : superpage_entries_2_valid_0; // @[TLB.scala 224:40]
  assign _GEN_471 = _T_1385 ? _GEN_371 : superpage_entries_3_valid_0; // @[TLB.scala 224:40]
  assign _GEN_473 = _T_1385 ? _GEN_373 : sectored_entries_0_valid_0; // @[TLB.scala 224:40]
  assign _GEN_474 = _T_1385 ? _GEN_374 : sectored_entries_0_valid_1; // @[TLB.scala 224:40]
  assign _GEN_475 = _T_1385 ? _GEN_375 : sectored_entries_0_valid_2; // @[TLB.scala 224:40]
  assign _GEN_476 = _T_1385 ? _GEN_376 : sectored_entries_0_valid_3; // @[TLB.scala 224:40]
  assign _GEN_483 = _T_1385 ? _GEN_383 : sectored_entries_1_valid_0; // @[TLB.scala 224:40]
  assign _GEN_484 = _T_1385 ? _GEN_384 : sectored_entries_1_valid_1; // @[TLB.scala 224:40]
  assign _GEN_485 = _T_1385 ? _GEN_385 : sectored_entries_1_valid_2; // @[TLB.scala 224:40]
  assign _GEN_486 = _T_1385 ? _GEN_386 : sectored_entries_1_valid_3; // @[TLB.scala 224:40]
  assign _GEN_493 = _T_1385 ? _GEN_393 : sectored_entries_2_valid_0; // @[TLB.scala 224:40]
  assign _GEN_494 = _T_1385 ? _GEN_394 : sectored_entries_2_valid_1; // @[TLB.scala 224:40]
  assign _GEN_495 = _T_1385 ? _GEN_395 : sectored_entries_2_valid_2; // @[TLB.scala 224:40]
  assign _GEN_496 = _T_1385 ? _GEN_396 : sectored_entries_2_valid_3; // @[TLB.scala 224:40]
  assign _GEN_503 = _T_1385 ? _GEN_403 : sectored_entries_3_valid_0; // @[TLB.scala 224:40]
  assign _GEN_504 = _T_1385 ? _GEN_404 : sectored_entries_3_valid_1; // @[TLB.scala 224:40]
  assign _GEN_505 = _T_1385 ? _GEN_405 : sectored_entries_3_valid_2; // @[TLB.scala 224:40]
  assign _GEN_506 = _T_1385 ? _GEN_406 : sectored_entries_3_valid_3; // @[TLB.scala 224:40]
  assign _GEN_513 = _T_1385 ? _GEN_413 : sectored_entries_4_valid_0; // @[TLB.scala 224:40]
  assign _GEN_514 = _T_1385 ? _GEN_414 : sectored_entries_4_valid_1; // @[TLB.scala 224:40]
  assign _GEN_515 = _T_1385 ? _GEN_415 : sectored_entries_4_valid_2; // @[TLB.scala 224:40]
  assign _GEN_516 = _T_1385 ? _GEN_416 : sectored_entries_4_valid_3; // @[TLB.scala 224:40]
  assign _GEN_523 = _T_1385 ? _GEN_423 : sectored_entries_5_valid_0; // @[TLB.scala 224:40]
  assign _GEN_524 = _T_1385 ? _GEN_424 : sectored_entries_5_valid_1; // @[TLB.scala 224:40]
  assign _GEN_525 = _T_1385 ? _GEN_425 : sectored_entries_5_valid_2; // @[TLB.scala 224:40]
  assign _GEN_526 = _T_1385 ? _GEN_426 : sectored_entries_5_valid_3; // @[TLB.scala 224:40]
  assign _GEN_533 = _T_1385 ? _GEN_433 : sectored_entries_6_valid_0; // @[TLB.scala 224:40]
  assign _GEN_534 = _T_1385 ? _GEN_434 : sectored_entries_6_valid_1; // @[TLB.scala 224:40]
  assign _GEN_535 = _T_1385 ? _GEN_435 : sectored_entries_6_valid_2; // @[TLB.scala 224:40]
  assign _GEN_536 = _T_1385 ? _GEN_436 : sectored_entries_6_valid_3; // @[TLB.scala 224:40]
  assign _GEN_543 = _T_1385 ? _GEN_443 : sectored_entries_7_valid_0; // @[TLB.scala 224:40]
  assign _GEN_544 = _T_1385 ? _GEN_444 : sectored_entries_7_valid_1; // @[TLB.scala 224:40]
  assign _GEN_545 = _T_1385 ? _GEN_445 : sectored_entries_7_valid_2; // @[TLB.scala 224:40]
  assign _GEN_546 = _T_1385 ? _GEN_446 : sectored_entries_7_valid_3; // @[TLB.scala 224:40]
  assign _T_2136 = {_GEN_55[11],_GEN_51[11],_GEN_47[11],_GEN_43[11],_GEN_39[11],_GEN_35[11]}; // @[Cat.scala 30:58]
  assign ptw_ae_array = {1'h0,special_entry_data_0[11],superpage_entries_3_data_0[11],superpage_entries_2_data_0[11],superpage_entries_1_data_0[11],superpage_entries_0_data_0[11],_GEN_63[11],_GEN_59[11],_T_2136}; // @[Cat.scala 30:58]
  assign _T_2150 = {_GEN_55[13],_GEN_51[13],_GEN_47[13],_GEN_43[13],_GEN_39[13],_GEN_35[13]}; // @[Cat.scala 30:58]
  assign _T_2157 = {special_entry_data_0[13],superpage_entries_3_data_0[13],superpage_entries_2_data_0[13],superpage_entries_1_data_0[13],superpage_entries_0_data_0[13],_GEN_63[13],_GEN_59[13],_T_2150}; // @[Cat.scala 30:58]
  assign priv_x_ok = priv_s ? ~_T_2157 : _T_2157; // @[TLB.scala 307:22]
  assign _T_2214 = {_GEN_55[9],_GEN_51[9],_GEN_47[9],_GEN_43[9],_GEN_39[9],_GEN_35[9]}; // @[Cat.scala 30:58]
  assign _T_2221 = {special_entry_data_0[9],superpage_entries_3_data_0[9],superpage_entries_2_data_0[9],superpage_entries_1_data_0[9],superpage_entries_0_data_0[9],_GEN_63[9],_GEN_59[9],_T_2214}; // @[Cat.scala 30:58]
  assign _T_2250 = priv_x_ok & _T_2221; // @[TLB.scala 310:39]
  assign x_array = {1'h1,_T_2250}; // @[Cat.scala 30:58]
  assign _T_2280 = prot_x ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign _T_2285 = {_GEN_55[6],_GEN_51[6],_GEN_47[6],_GEN_43[6],_GEN_39[6],_GEN_35[6]}; // @[Cat.scala 30:58]
  assign _T_2292 = {_T_2280,superpage_entries_3_data_0[6],superpage_entries_2_data_0[6],superpage_entries_1_data_0[6],superpage_entries_0_data_0[6],_GEN_63[6],_GEN_59[6],_T_2285}; // @[Cat.scala 30:58]
  assign px_array = _T_2292 | ptw_ae_array; // @[TLB.scala 313:87]
  assign _T_2333 = cacheable ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign _T_2338 = {_GEN_55[1],_GEN_51[1],_GEN_47[1],_GEN_43[1],_GEN_39[1],_GEN_35[1]}; // @[Cat.scala 30:58]
  assign c_array = {_T_2333,superpage_entries_3_data_0[1],superpage_entries_2_data_0[1],superpage_entries_1_data_0[1],superpage_entries_0_data_0[1],_GEN_63[1],_GEN_59[1],_T_2338}; // @[Cat.scala 30:58]
  assign _T_2364 = $signed(io_req_bits_vaddr) < 40'sh0; // @[TLB.scala 323:37]
  assign _T_2365 = io_req_bits_vaddr[38:12]; // @[TLB.scala 323:53]
  assign _T_2366 = $signed(_T_2365) < 27'sh0; // @[TLB.scala 323:60]
  assign _T_2367 = _T_2364 != _T_2366; // @[TLB.scala 323:44]
  assign bad_va = vm_enabled & _T_2367; // @[TLB.scala 321:27]
  assign _T_2549 = x_array | ptw_ae_array; // @[TLB.scala 338:33]
  assign pf_inst_array = ~_T_2549; // @[TLB.scala 338:23]
  assign tlb_hit = real_hits != 13'h0; // @[TLB.scala 340:27]
  assign _T_2551 = vm_enabled & ~bad_va; // @[TLB.scala 341:29]
  assign tlb_miss = _T_2551 & ~tlb_hit; // @[TLB.scala 341:40]
  assign _T_2557 = io_req_valid & vm_enabled; // @[TLB.scala 345:22]
  assign _T_2558 = sector_hits_0 | sector_hits_1; // @[package.scala 63:59]
  assign _T_2559 = _T_2558 | sector_hits_2; // @[package.scala 63:59]
  assign _T_2560 = _T_2559 | sector_hits_3; // @[package.scala 63:59]
  assign _T_2561 = _T_2560 | sector_hits_4; // @[package.scala 63:59]
  assign _T_2562 = _T_2561 | sector_hits_5; // @[package.scala 63:59]
  assign _T_2563 = _T_2562 | sector_hits_6; // @[package.scala 63:59]
  assign _T_2564 = _T_2563 | sector_hits_7; // @[package.scala 63:59]
  assign _T_2571 = {sector_hits_7,sector_hits_6,sector_hits_5,sector_hits_4,sector_hits_3,sector_hits_2,sector_hits_1,sector_hits_0}; // @[Cat.scala 30:58]
  assign _T_2574 = _T_2571[7:4] != 4'h0; // @[OneHot.scala 28:14]
  assign _T_2575 = _T_2571[7:4] | _T_2571[3:0]; // @[OneHot.scala 28:28]
  assign _T_2578 = _T_2575[3:2] != 2'h0; // @[OneHot.scala 28:14]
  assign _T_2579 = _T_2575[3:2] | _T_2575[1:0]; // @[OneHot.scala 28:28]
  assign _T_2582 = {_T_2574,_T_2578,_T_2579[1]}; // @[Cat.scala 30:58]
  assign _T_2583 = {_T_2554, 1'h0}; // @[Replacement.scala 46:28]
  assign _T_2587 = _T_2583 | 8'h2; // @[Replacement.scala 50:37]
  assign _T_2589 = ~_T_2583 | 8'h2; // @[Replacement.scala 50:37]
  assign _T_2591 = _T_2582[2] ? ~_T_2589 : _T_2587; // @[Replacement.scala 50:37]
  assign _T_2592 = {1'h1,_T_2582[2]}; // @[Cat.scala 30:58]
  assign _T_2595 = 4'h1 << _T_2592; // @[Replacement.scala 50:37]
  assign _GEN_1001 = {{4'd0}, _T_2595}; // @[Replacement.scala 50:37]
  assign _T_2596 = _T_2591 | _GEN_1001; // @[Replacement.scala 50:37]
  assign _T_2598 = ~_T_2591 | _GEN_1001; // @[Replacement.scala 50:37]
  assign _T_2600 = _T_2582[1] ? ~_T_2598 : _T_2596; // @[Replacement.scala 50:37]
  assign _T_2601 = {1'h1,_T_2582[2],_T_2582[1]}; // @[Cat.scala 30:58]
  assign _T_2604 = 8'h1 << _T_2601; // @[Replacement.scala 50:37]
  assign _T_2605 = _T_2600 | _T_2604; // @[Replacement.scala 50:37]
  assign _T_2607 = ~_T_2600 | _T_2604; // @[Replacement.scala 50:37]
  assign _T_2609 = _T_2582[0] ? ~_T_2607 : _T_2605; // @[Replacement.scala 50:37]
  assign _T_2612 = superpage_hits_0 | superpage_hits_1; // @[package.scala 63:59]
  assign _T_2613 = _T_2612 | superpage_hits_2; // @[package.scala 63:59]
  assign _T_2614 = _T_2613 | superpage_hits_3; // @[package.scala 63:59]
  assign _T_2617 = {superpage_hits_3,superpage_hits_2,superpage_hits_1,superpage_hits_0}; // @[Cat.scala 30:58]
  assign _T_2620 = _T_2617[3:2] != 2'h0; // @[OneHot.scala 28:14]
  assign _T_2621 = _T_2617[3:2] | _T_2617[1:0]; // @[OneHot.scala 28:28]
  assign _T_2623 = {_T_2620,_T_2621[1]}; // @[Cat.scala 30:58]
  assign _T_2624 = {_T_2556, 1'h0}; // @[Replacement.scala 46:28]
  assign _T_2628 = _T_2624 | 4'h2; // @[Replacement.scala 50:37]
  assign _T_2630 = ~_T_2624 | 4'h2; // @[Replacement.scala 50:37]
  assign _T_2632 = _T_2623[1] ? ~_T_2630 : _T_2628; // @[Replacement.scala 50:37]
  assign _T_2633 = {1'h1,_T_2623[1]}; // @[Cat.scala 30:58]
  assign _T_2636 = 4'h1 << _T_2633; // @[Replacement.scala 50:37]
  assign _T_2637 = _T_2632 | _T_2636; // @[Replacement.scala 50:37]
  assign _T_2639 = ~_T_2632 | _T_2636; // @[Replacement.scala 50:37]
  assign _T_2641 = _T_2623[0] ? ~_T_2639 : _T_2637; // @[Replacement.scala 50:37]
  assign _T_2653 = real_hits[1] | real_hits[2]; // @[Misc.scala 187:16]
  assign _T_2655 = real_hits[1] & real_hits[2]; // @[Misc.scala 187:61]
  assign _T_2657 = real_hits[0] | _T_2653; // @[Misc.scala 187:16]
  assign _T_2659 = real_hits[0] & _T_2653; // @[Misc.scala 187:61]
  assign _T_2660 = _T_2655 | _T_2659; // @[Misc.scala 187:49]
  assign _T_2669 = real_hits[4] | real_hits[5]; // @[Misc.scala 187:16]
  assign _T_2671 = real_hits[4] & real_hits[5]; // @[Misc.scala 187:61]
  assign _T_2673 = real_hits[3] | _T_2669; // @[Misc.scala 187:16]
  assign _T_2675 = real_hits[3] & _T_2669; // @[Misc.scala 187:61]
  assign _T_2676 = _T_2671 | _T_2675; // @[Misc.scala 187:49]
  assign _T_2677 = _T_2657 | _T_2673; // @[Misc.scala 187:16]
  assign _T_2678 = _T_2660 | _T_2676; // @[Misc.scala 187:37]
  assign _T_2679 = _T_2657 & _T_2673; // @[Misc.scala 187:61]
  assign _T_2680 = _T_2678 | _T_2679; // @[Misc.scala 187:49]
  assign _T_2690 = real_hits[7] | real_hits[8]; // @[Misc.scala 187:16]
  assign _T_2692 = real_hits[7] & real_hits[8]; // @[Misc.scala 187:61]
  assign _T_2694 = real_hits[6] | _T_2690; // @[Misc.scala 187:16]
  assign _T_2696 = real_hits[6] & _T_2690; // @[Misc.scala 187:61]
  assign _T_2697 = _T_2692 | _T_2696; // @[Misc.scala 187:49]
  assign _T_2704 = real_hits[9] | real_hits[10]; // @[Misc.scala 187:16]
  assign _T_2706 = real_hits[9] & real_hits[10]; // @[Misc.scala 187:61]
  assign _T_2713 = real_hits[11] | real_hits[12]; // @[Misc.scala 187:16]
  assign _T_2715 = real_hits[11] & real_hits[12]; // @[Misc.scala 187:61]
  assign _T_2717 = _T_2704 | _T_2713; // @[Misc.scala 187:16]
  assign _T_2718 = _T_2706 | _T_2715; // @[Misc.scala 187:37]
  assign _T_2719 = _T_2704 & _T_2713; // @[Misc.scala 187:61]
  assign _T_2720 = _T_2718 | _T_2719; // @[Misc.scala 187:49]
  assign _T_2721 = _T_2694 | _T_2717; // @[Misc.scala 187:16]
  assign _T_2722 = _T_2697 | _T_2720; // @[Misc.scala 187:37]
  assign _T_2723 = _T_2694 & _T_2717; // @[Misc.scala 187:61]
  assign _T_2724 = _T_2722 | _T_2723; // @[Misc.scala 187:49]
  assign _T_2726 = _T_2680 | _T_2724; // @[Misc.scala 187:37]
  assign _T_2727 = _T_2677 & _T_2721; // @[Misc.scala 187:61]
  assign multipleHits = _T_2726 | _T_2727; // @[Misc.scala 187:49]
  assign _T_2783 = pf_inst_array & hits; // @[TLB.scala 360:47]
  assign _T_2784 = _T_2783 != 14'h0; // @[TLB.scala 360:55]
  assign _T_2791 = ~px_array & hits; // @[TLB.scala 363:33]
  assign _T_2797 = c_array & hits; // @[TLB.scala 367:33]
  assign _T_2802 = io_ptw_resp_valid | tlb_miss; // @[TLB.scala 369:29]
  assign _T_2808 = io_req_ready & io_req_valid; // @[Decoupled.scala 37:37]
  assign _T_2809 = _T_2808 & tlb_miss; // @[TLB.scala 385:25]
  assign _T_2814 = {{1'd0}, _T_2624[3:1]}; // @[Replacement.scala 61:48]
  assign _T_2817 = {1'h1,_T_2814[0]}; // @[Cat.scala 30:58]
  assign _T_2821 = _T_2624 >> _T_2817; // @[Replacement.scala 61:48]
  assign _T_2824 = {1'h1,_T_2814[0],_T_2821[0]}; // @[Cat.scala 30:58]
  assign _T_2828 = {superpage_entries_3_valid_0,superpage_entries_2_valid_0,superpage_entries_1_valid_0,superpage_entries_0_valid_0}; // @[Cat.scala 30:58]
  assign _T_2830 = ~_T_2828 == 4'h0; // @[TLB.scala 440:16]
  assign _T_2832 = ~_T_2828[0]; // @[OneHot.scala 39:40]
  assign _T_2833 = ~_T_2828[1]; // @[OneHot.scala 39:40]
  assign _T_2834 = ~_T_2828[2]; // @[OneHot.scala 39:40]
  assign _T_2844 = {{1'd0}, _T_2583[7:1]}; // @[Replacement.scala 61:48]
  assign _T_2847 = {1'h1,_T_2844[0]}; // @[Cat.scala 30:58]
  assign _T_2851 = _T_2583 >> _T_2847; // @[Replacement.scala 61:48]
  assign _T_2854 = {1'h1,_T_2844[0],_T_2851[0]}; // @[Cat.scala 30:58]
  assign _T_2858 = _T_2583 >> _T_2854; // @[Replacement.scala 61:48]
  assign _T_2861 = {1'h1,_T_2844[0],_T_2851[0],_T_2858[0]}; // @[Cat.scala 30:58]
  assign _T_2893 = {_T_766,_T_760,_T_754,_T_748,_T_742,_T_736,_T_730,_T_724}; // @[Cat.scala 30:58]
  assign _T_2895 = ~_T_2893 == 8'h0; // @[TLB.scala 440:16]
  assign _T_2897 = ~_T_2893[0]; // @[OneHot.scala 39:40]
  assign _T_2898 = ~_T_2893[1]; // @[OneHot.scala 39:40]
  assign _T_2899 = ~_T_2893[2]; // @[OneHot.scala 39:40]
  assign _T_2900 = ~_T_2893[3]; // @[OneHot.scala 39:40]
  assign _T_2901 = ~_T_2893[4]; // @[OneHot.scala 39:40]
  assign _T_2902 = ~_T_2893[5]; // @[OneHot.scala 39:40]
  assign _T_2903 = ~_T_2893[6]; // @[OneHot.scala 39:40]
  assign _T_2940 = state == 2'h2; // @[TLB.scala 399:17]
  assign _T_2941 = _T_2940 & io_sfence_valid; // @[TLB.scala 399:28]
  assign _T_2946 = io_sfence_bits_addr[38:12] == vpn; // @[TLB.scala 414:72]
  assign _T_2947 = ~io_sfence_bits_rs1 | _T_2946; // @[TLB.scala 414:34]
  assign _T_2949 = _T_2947 | reset; // @[TLB.scala 414:13]
  assign _T_2957 = _T_725[26:18] == 9'h0; // @[TLB.scala 150:63]
  assign _GEN_652 = sectored_entries_0_data_0[12] ? _GEN_473 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_653 = sectored_entries_0_data_1[12] ? _GEN_474 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_654 = sectored_entries_0_data_2[12] ? _GEN_475 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_655 = sectored_entries_0_data_3[12] ? _GEN_476 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_656 = io_sfence_bits_rs2 & _GEN_652; // @[TLB.scala 417:40]
  assign _GEN_657 = io_sfence_bits_rs2 & _GEN_653; // @[TLB.scala 417:40]
  assign _GEN_658 = io_sfence_bits_rs2 & _GEN_654; // @[TLB.scala 417:40]
  assign _GEN_659 = io_sfence_bits_rs2 & _GEN_655; // @[TLB.scala 417:40]
  assign _T_3128 = _T_731[26:18] == 9'h0; // @[TLB.scala 150:63]
  assign _GEN_680 = sectored_entries_1_data_0[12] ? _GEN_483 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_681 = sectored_entries_1_data_1[12] ? _GEN_484 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_682 = sectored_entries_1_data_2[12] ? _GEN_485 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_683 = sectored_entries_1_data_3[12] ? _GEN_486 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_684 = io_sfence_bits_rs2 & _GEN_680; // @[TLB.scala 417:40]
  assign _GEN_685 = io_sfence_bits_rs2 & _GEN_681; // @[TLB.scala 417:40]
  assign _GEN_686 = io_sfence_bits_rs2 & _GEN_682; // @[TLB.scala 417:40]
  assign _GEN_687 = io_sfence_bits_rs2 & _GEN_683; // @[TLB.scala 417:40]
  assign _T_3299 = _T_737[26:18] == 9'h0; // @[TLB.scala 150:63]
  assign _GEN_708 = sectored_entries_2_data_0[12] ? _GEN_493 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_709 = sectored_entries_2_data_1[12] ? _GEN_494 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_710 = sectored_entries_2_data_2[12] ? _GEN_495 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_711 = sectored_entries_2_data_3[12] ? _GEN_496 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_712 = io_sfence_bits_rs2 & _GEN_708; // @[TLB.scala 417:40]
  assign _GEN_713 = io_sfence_bits_rs2 & _GEN_709; // @[TLB.scala 417:40]
  assign _GEN_714 = io_sfence_bits_rs2 & _GEN_710; // @[TLB.scala 417:40]
  assign _GEN_715 = io_sfence_bits_rs2 & _GEN_711; // @[TLB.scala 417:40]
  assign _T_3470 = _T_743[26:18] == 9'h0; // @[TLB.scala 150:63]
  assign _GEN_736 = sectored_entries_3_data_0[12] ? _GEN_503 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_737 = sectored_entries_3_data_1[12] ? _GEN_504 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_738 = sectored_entries_3_data_2[12] ? _GEN_505 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_739 = sectored_entries_3_data_3[12] ? _GEN_506 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_740 = io_sfence_bits_rs2 & _GEN_736; // @[TLB.scala 417:40]
  assign _GEN_741 = io_sfence_bits_rs2 & _GEN_737; // @[TLB.scala 417:40]
  assign _GEN_742 = io_sfence_bits_rs2 & _GEN_738; // @[TLB.scala 417:40]
  assign _GEN_743 = io_sfence_bits_rs2 & _GEN_739; // @[TLB.scala 417:40]
  assign _T_3641 = _T_749[26:18] == 9'h0; // @[TLB.scala 150:63]
  assign _GEN_764 = sectored_entries_4_data_0[12] ? _GEN_513 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_765 = sectored_entries_4_data_1[12] ? _GEN_514 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_766 = sectored_entries_4_data_2[12] ? _GEN_515 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_767 = sectored_entries_4_data_3[12] ? _GEN_516 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_768 = io_sfence_bits_rs2 & _GEN_764; // @[TLB.scala 417:40]
  assign _GEN_769 = io_sfence_bits_rs2 & _GEN_765; // @[TLB.scala 417:40]
  assign _GEN_770 = io_sfence_bits_rs2 & _GEN_766; // @[TLB.scala 417:40]
  assign _GEN_771 = io_sfence_bits_rs2 & _GEN_767; // @[TLB.scala 417:40]
  assign _T_3812 = _T_755[26:18] == 9'h0; // @[TLB.scala 150:63]
  assign _GEN_792 = sectored_entries_5_data_0[12] ? _GEN_523 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_793 = sectored_entries_5_data_1[12] ? _GEN_524 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_794 = sectored_entries_5_data_2[12] ? _GEN_525 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_795 = sectored_entries_5_data_3[12] ? _GEN_526 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_796 = io_sfence_bits_rs2 & _GEN_792; // @[TLB.scala 417:40]
  assign _GEN_797 = io_sfence_bits_rs2 & _GEN_793; // @[TLB.scala 417:40]
  assign _GEN_798 = io_sfence_bits_rs2 & _GEN_794; // @[TLB.scala 417:40]
  assign _GEN_799 = io_sfence_bits_rs2 & _GEN_795; // @[TLB.scala 417:40]
  assign _T_3983 = _T_761[26:18] == 9'h0; // @[TLB.scala 150:63]
  assign _GEN_820 = sectored_entries_6_data_0[12] ? _GEN_533 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_821 = sectored_entries_6_data_1[12] ? _GEN_534 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_822 = sectored_entries_6_data_2[12] ? _GEN_535 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_823 = sectored_entries_6_data_3[12] ? _GEN_536 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_824 = io_sfence_bits_rs2 & _GEN_820; // @[TLB.scala 417:40]
  assign _GEN_825 = io_sfence_bits_rs2 & _GEN_821; // @[TLB.scala 417:40]
  assign _GEN_826 = io_sfence_bits_rs2 & _GEN_822; // @[TLB.scala 417:40]
  assign _GEN_827 = io_sfence_bits_rs2 & _GEN_823; // @[TLB.scala 417:40]
  assign _T_4154 = _T_767[26:18] == 9'h0; // @[TLB.scala 150:63]
  assign _GEN_848 = sectored_entries_7_data_0[12] ? _GEN_543 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_849 = sectored_entries_7_data_1[12] ? _GEN_544 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_850 = sectored_entries_7_data_2[12] ? _GEN_545 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_851 = sectored_entries_7_data_3[12] ? _GEN_546 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_852 = io_sfence_bits_rs2 & _GEN_848; // @[TLB.scala 417:40]
  assign _GEN_853 = io_sfence_bits_rs2 & _GEN_849; // @[TLB.scala 417:40]
  assign _GEN_854 = io_sfence_bits_rs2 & _GEN_850; // @[TLB.scala 417:40]
  assign _GEN_855 = io_sfence_bits_rs2 & _GEN_851; // @[TLB.scala 417:40]
  assign _GEN_861 = superpage_entries_0_data_0[12] ? _GEN_459 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_862 = io_sfence_bits_rs2 & _GEN_861; // @[TLB.scala 417:40]
  assign _GEN_865 = superpage_entries_1_data_0[12] ? _GEN_463 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_866 = io_sfence_bits_rs2 & _GEN_865; // @[TLB.scala 417:40]
  assign _GEN_869 = superpage_entries_2_data_0[12] ? _GEN_467 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_870 = io_sfence_bits_rs2 & _GEN_869; // @[TLB.scala 417:40]
  assign _GEN_873 = superpage_entries_3_data_0[12] ? _GEN_471 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_874 = io_sfence_bits_rs2 & _GEN_873; // @[TLB.scala 417:40]
  assign _GEN_877 = special_entry_data_0[12] ? _GEN_455 : 1'h0; // @[TLB.scala 158:21]
  assign _GEN_878 = io_sfence_bits_rs2 & _GEN_877; // @[TLB.scala 417:40]
  assign _T_4530 = multipleHits | reset; // @[TLB.scala 421:24]
  assign io_req_ready = state == 2'h0; // @[TLB.scala 357:16]
  assign io_resp_miss = _T_2802 | multipleHits; // @[TLB.scala 369:16]
  assign io_resp_paddr = {ppn,io_req_bits_vaddr[11:0]}; // @[TLB.scala 370:17]
  assign io_resp_pf_inst = bad_va | _T_2784; // @[TLB.scala 360:19]
  assign io_resp_ae_inst = _T_2791 != 14'h0; // @[TLB.scala 363:19]
  assign io_resp_cacheable = _T_2797 != 14'h0; // @[TLB.scala 367:21]
  assign io_ptw_req_valid = state == 2'h1; // @[TLB.scala 372:20]
  assign io_ptw_req_bits_valid = ~io_kill; // @[TLB.scala 373:25]
  assign io_ptw_req_bits_bits_addr = r_refill_tag; // @[TLB.scala 374:29]
  assign pmp_io_prv = io_ptw_resp_valid ? 2'h1 : io_ptw_status_prv; // @[TLB.scala 194:14]
  assign pmp_io_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_addr = io_ptw_pmp_0_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_mask = io_ptw_pmp_0_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_addr = io_ptw_pmp_1_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_mask = io_ptw_pmp_1_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_addr = io_ptw_pmp_2_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_mask = io_ptw_pmp_2_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_addr = io_ptw_pmp_3_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_mask = io_ptw_pmp_3_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_addr = io_ptw_pmp_4_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_mask = io_ptw_pmp_4_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_addr = io_ptw_pmp_5_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_mask = io_ptw_pmp_5_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_addr = io_ptw_pmp_6_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_mask = io_ptw_pmp_6_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_addr = io_ptw_pmp_7_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_mask = io_ptw_pmp_7_mask; // @[TLB.scala 193:14]
  assign pmp_io_addr = mpu_physaddr[31:0]; // @[TLB.scala 191:15]
  assign TLB_1_cov_read_addr = TLB_1_state;
  assign TLB_1_cov_read_data = TLB_1_cov[TLB_1_cov_read_addr]; // @[Coverage map for TLB_1]
  assign TLB_1_cov_write_data = 1'h1;
  assign TLB_1_cov_write_addr = TLB_1_state;
  assign TLB_1_cov_write_mask = 1'h1;
  assign TLB_1_cov_write_en = 1'h1;
  assign mux_cond_0 = sectored_entries_0_data_0[0];
  assign mux_cond_1 = ~sectored_entries_3_data_3[12];
  assign mux_cond_2 = sectored_entries_1_data_0[0];
  assign mux_cond_3 = ~sectored_entries_4_data_3[12];
  assign mux_cond_4 = ~superpage_entries_0_data_0[12];
  assign mux_cond_5 = ~sectored_entries_2_data_1[12];
  assign mux_cond_6 = sectored_entries_2_data_3[0];
  assign mux_cond_7 = ~sectored_entries_4_data_2[12];
  assign mux_cond_8 = ~sectored_entries_5_data_1[12];
  assign mux_cond_9 = sectored_entries_0_data_1[0];
  assign mux_cond_10 = sectored_entries_3_data_1[0];
  assign mux_cond_11 = ~sectored_entries_4_data_1[12];
  assign mux_cond_12 = sectored_entries_7_data_1[0];
  assign mux_cond_13 = ~sectored_entries_0_data_3[12];
  assign mux_cond_14 = ~sectored_entries_1_data_2[12];
  assign mux_cond_15 = sectored_entries_5_data_2[0];
  assign mux_cond_16 = ~special_entry_data_0[12];
  assign mux_cond_17 = sectored_entries_5_data_3[0];
  assign mux_cond_18 = sectored_entries_6_data_1[0];
  assign mux_cond_19 = ~sectored_entries_2_data_3[12];
  assign mux_cond_20 = ~superpage_entries_1_data_0[12];
  assign mux_cond_21 = ~sectored_entries_3_data_0[12];
  assign mux_cond_22 = sectored_entries_4_data_0[0];
  assign mux_cond_23 = sectored_entries_7_data_3[0];
  assign mux_cond_24 = ~sectored_entries_1_data_1[12];
  assign mux_cond_25 = sectored_entries_2_data_0[0];
  assign mux_cond_26 = ~sectored_entries_1_data_0[12];
  assign mux_cond_27 = sectored_entries_1_data_2[0];
  assign mux_cond_28 = ~sectored_entries_5_data_2[12];
  assign mux_cond_29 = sectored_entries_3_data_2[0];
  assign mux_cond_30 = ~sectored_entries_3_data_2[12];
  assign mux_cond_31 = ~sectored_entries_7_data_2[12];
  assign mux_cond_32 = ~sectored_entries_2_data_2[12];
  assign mux_cond_33 = sectored_entries_4_data_3[0];
  assign mux_cond_34 = sectored_entries_5_data_0[0];
  assign mux_cond_35 = sectored_entries_7_data_0[0];
  assign mux_cond_36 = sectored_entries_2_data_2[0];
  assign mux_cond_37 = sectored_entries_6_data_3[0];
  assign mux_cond_38 = prot_x;
  assign mux_cond_39 = ~superpage_entries_3_data_0[12];
  assign mux_cond_40 = ~sectored_entries_7_data_3[12];
  assign mux_cond_41 = ~sectored_entries_7_data_1[12];
  assign mux_cond_42 = sectored_entries_1_data_1[0];
  assign mux_cond_43 = sectored_entries_0_data_3[0];
  assign mux_cond_44 = cacheable;
  assign mux_cond_45 = sectored_entries_5_data_1[0];
  assign mux_cond_46 = ~sectored_entries_5_data_3[12];
  assign mux_cond_47 = ~sectored_entries_0_data_2[12];
  assign mux_cond_48 = ~sectored_entries_1_data_3[12];
  assign mux_cond_49 = sectored_entries_6_data_2[0];
  assign mux_cond_50 = ~sectored_entries_4_data_0[12];
  assign mux_cond_51 = ~sectored_entries_0_data_0[12];
  assign mux_cond_52 = ~sectored_entries_7_data_0[12];
  assign mux_cond_53 = ~sectored_entries_3_data_1[12];
  assign mux_cond_54 = ~sectored_entries_5_data_0[12];
  assign mux_cond_55 = sectored_entries_3_data_0[0];
  assign mux_cond_56 = sectored_entries_7_data_2[0];
  assign mux_cond_57 = ~sectored_entries_2_data_0[12];
  assign mux_cond_58 = sectored_entries_4_data_2[0];
  assign mux_cond_59 = sectored_entries_1_data_3[0];
  assign mux_cond_60 = ~sectored_entries_6_data_2[12];
  assign mux_cond_61 = ~sectored_entries_6_data_0[12];
  assign mux_cond_62 = ~sectored_entries_0_data_1[12];
  assign mux_cond_63 = sectored_entries_3_data_3[0];
  assign mux_cond_64 = ~superpage_entries_2_data_0[12];
  assign mux_cond_65 = sectored_entries_6_data_0[0];
  assign mux_cond_66 = sectored_entries_4_data_1[0];
  assign mux_cond_67 = ~sectored_entries_6_data_3[12];
  assign mux_cond_68 = sectored_entries_0_data_2[0];
  assign mux_cond_69 = sectored_entries_2_data_1[0];
  assign mux_cond_70 = ~sectored_entries_6_data_1[12];
  assign r_superpage_repl_addr_shl = {r_superpage_repl_addr, 18'h0};
  assign r_superpage_repl_addr_pad = r_superpage_repl_addr_shl;
  assign state_shl = {state, 3'h0};
  assign state_pad = {15'h0,state_shl};
  assign r_sectored_repl_addr_shl = {r_sectored_repl_addr, 14'h0};
  assign r_sectored_repl_addr_pad = {3'h0,r_sectored_repl_addr_shl};
  assign r_sectored_hit_addr_shl = {r_sectored_hit_addr, 3'h0};
  assign r_sectored_hit_addr_pad = {14'h0,r_sectored_hit_addr_shl};
  assign special_entry_valid_0_shl = {special_entry_valid_0, 9'h0};
  assign special_entry_valid_0_pad = {10'h0,special_entry_valid_0_shl};
  assign special_entry_level_shl = {special_entry_level, 1'h0};
  assign special_entry_level_pad = {17'h0,special_entry_level_shl};
  assign r_sectored_hit_shl = {r_sectored_hit, 1'h0};
  assign r_sectored_hit_pad = {18'h0,r_sectored_hit_shl};
  assign mux_cond_0_shl = {mux_cond_0, 1'h0};
  assign mux_cond_0_pad = {18'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 3'h0};
  assign mux_cond_1_pad = {16'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 6'h0};
  assign mux_cond_2_pad = {13'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 14'h0};
  assign mux_cond_3_pad = {5'h0,mux_cond_3_shl};
  assign mux_cond_4_shl = {mux_cond_4, 17'h0};
  assign mux_cond_4_pad = {2'h0,mux_cond_4_shl};
  assign mux_cond_5_shl = {mux_cond_5, 19'h0};
  assign mux_cond_5_pad = mux_cond_5_shl;
  assign mux_cond_6_shl = {mux_cond_6, 7'h0};
  assign mux_cond_6_pad = {12'h0,mux_cond_6_shl};
  assign mux_cond_7_shl = {mux_cond_7, 16'h0};
  assign mux_cond_7_pad = {3'h0,mux_cond_7_shl};
  assign mux_cond_8_shl = {mux_cond_8, 7'h0};
  assign mux_cond_8_pad = {12'h0,mux_cond_8_shl};
  assign mux_cond_9_shl = {mux_cond_9, 10'h0};
  assign mux_cond_9_pad = {9'h0,mux_cond_9_shl};
  assign mux_cond_10_shl = {mux_cond_10, 14'h0};
  assign mux_cond_10_pad = {5'h0,mux_cond_10_shl};
  assign mux_cond_11_shl = {mux_cond_11, 9'h0};
  assign mux_cond_11_pad = {10'h0,mux_cond_11_shl};
  assign mux_cond_12_shl = {mux_cond_12, 9'h0};
  assign mux_cond_12_pad = {10'h0,mux_cond_12_shl};
  assign mux_cond_13_shl = {mux_cond_13, 9'h0};
  assign mux_cond_13_pad = {10'h0,mux_cond_13_shl};
  assign mux_cond_14_shl = {mux_cond_14, 14'h0};
  assign mux_cond_14_pad = {5'h0,mux_cond_14_shl};
  assign mux_cond_15_shl = {mux_cond_15, 8'h0};
  assign mux_cond_15_pad = {11'h0,mux_cond_15_shl};
  assign mux_cond_16_shl = {mux_cond_16, 15'h0};
  assign mux_cond_16_pad = {4'h0,mux_cond_16_shl};
  assign mux_cond_17_shl = {mux_cond_17, 10'h0};
  assign mux_cond_17_pad = {9'h0,mux_cond_17_shl};
  assign mux_cond_18_shl = mux_cond_18;
  assign mux_cond_18_pad = {19'h0,mux_cond_18_shl};
  assign mux_cond_19_shl = {mux_cond_19, 13'h0};
  assign mux_cond_19_pad = {6'h0,mux_cond_19_shl};
  assign mux_cond_20_shl = {mux_cond_20, 9'h0};
  assign mux_cond_20_pad = {10'h0,mux_cond_20_shl};
  assign mux_cond_21_shl = {mux_cond_21, 16'h0};
  assign mux_cond_21_pad = {3'h0,mux_cond_21_shl};
  assign mux_cond_22_shl = {mux_cond_22, 5'h0};
  assign mux_cond_22_pad = {14'h0,mux_cond_22_shl};
  assign mux_cond_23_shl = {mux_cond_23, 19'h0};
  assign mux_cond_23_pad = mux_cond_23_shl;
  assign mux_cond_24_shl = {mux_cond_24, 1'h0};
  assign mux_cond_24_pad = {18'h0,mux_cond_24_shl};
  assign mux_cond_25_shl = {mux_cond_25, 8'h0};
  assign mux_cond_25_pad = {11'h0,mux_cond_25_shl};
  assign mux_cond_26_shl = {mux_cond_26, 12'h0};
  assign mux_cond_26_pad = {7'h0,mux_cond_26_shl};
  assign mux_cond_27_shl = {mux_cond_27, 14'h0};
  assign mux_cond_27_pad = {5'h0,mux_cond_27_shl};
  assign mux_cond_28_shl = {mux_cond_28, 7'h0};
  assign mux_cond_28_pad = {12'h0,mux_cond_28_shl};
  assign mux_cond_29_shl = {mux_cond_29, 11'h0};
  assign mux_cond_29_pad = {8'h0,mux_cond_29_shl};
  assign mux_cond_30_shl = {mux_cond_30, 8'h0};
  assign mux_cond_30_pad = {11'h0,mux_cond_30_shl};
  assign mux_cond_31_shl = {mux_cond_31, 6'h0};
  assign mux_cond_31_pad = {13'h0,mux_cond_31_shl};
  assign mux_cond_32_shl = {mux_cond_32, 6'h0};
  assign mux_cond_32_pad = {13'h0,mux_cond_32_shl};
  assign mux_cond_33_shl = {mux_cond_33, 6'h0};
  assign mux_cond_33_pad = {13'h0,mux_cond_33_shl};
  assign mux_cond_34_shl = {mux_cond_34, 16'h0};
  assign mux_cond_34_pad = {3'h0,mux_cond_34_shl};
  assign mux_cond_35_shl = {mux_cond_35, 11'h0};
  assign mux_cond_35_pad = {8'h0,mux_cond_35_shl};
  assign mux_cond_36_shl = {mux_cond_36, 4'h0};
  assign mux_cond_36_pad = {15'h0,mux_cond_36_shl};
  assign mux_cond_37_shl = {mux_cond_37, 7'h0};
  assign mux_cond_37_pad = {12'h0,mux_cond_37_shl};
  assign mux_cond_38_shl = {mux_cond_38, 11'h0};
  assign mux_cond_38_pad = {8'h0,mux_cond_38_shl};
  assign mux_cond_39_shl = {mux_cond_39, 14'h0};
  assign mux_cond_39_pad = {5'h0,mux_cond_39_shl};
  assign mux_cond_40_shl = {mux_cond_40, 7'h0};
  assign mux_cond_40_pad = {12'h0,mux_cond_40_shl};
  assign mux_cond_41_shl = {mux_cond_41, 9'h0};
  assign mux_cond_41_pad = {10'h0,mux_cond_41_shl};
  assign mux_cond_42_shl = {mux_cond_42, 1'h0};
  assign mux_cond_42_pad = {18'h0,mux_cond_42_shl};
  assign mux_cond_43_shl = {mux_cond_43, 4'h0};
  assign mux_cond_43_pad = {15'h0,mux_cond_43_shl};
  assign mux_cond_44_shl = {mux_cond_44, 6'h0};
  assign mux_cond_44_pad = {13'h0,mux_cond_44_shl};
  assign mux_cond_45_shl = {mux_cond_45, 15'h0};
  assign mux_cond_45_pad = {4'h0,mux_cond_45_shl};
  assign mux_cond_46_shl = {mux_cond_46, 18'h0};
  assign mux_cond_46_pad = {1'h0,mux_cond_46_shl};
  assign mux_cond_47_shl = {mux_cond_47, 2'h0};
  assign mux_cond_47_pad = {17'h0,mux_cond_47_shl};
  assign mux_cond_48_shl = {mux_cond_48, 11'h0};
  assign mux_cond_48_pad = {8'h0,mux_cond_48_shl};
  assign mux_cond_49_shl = {mux_cond_49, 14'h0};
  assign mux_cond_49_pad = {5'h0,mux_cond_49_shl};
  assign mux_cond_50_shl = {mux_cond_50, 15'h0};
  assign mux_cond_50_pad = {4'h0,mux_cond_50_shl};
  assign mux_cond_51_shl = {mux_cond_51, 9'h0};
  assign mux_cond_51_pad = {10'h0,mux_cond_51_shl};
  assign mux_cond_52_shl = {mux_cond_52, 18'h0};
  assign mux_cond_52_pad = {1'h0,mux_cond_52_shl};
  assign mux_cond_53_shl = {mux_cond_53, 18'h0};
  assign mux_cond_53_pad = {1'h0,mux_cond_53_shl};
  assign mux_cond_54_shl = {mux_cond_54, 10'h0};
  assign mux_cond_54_pad = {9'h0,mux_cond_54_shl};
  assign mux_cond_55_shl = {mux_cond_55, 9'h0};
  assign mux_cond_55_pad = {10'h0,mux_cond_55_shl};
  assign mux_cond_56_shl = mux_cond_56;
  assign mux_cond_56_pad = {19'h0,mux_cond_56_shl};
  assign mux_cond_57_shl = {mux_cond_57, 3'h0};
  assign mux_cond_57_pad = {16'h0,mux_cond_57_shl};
  assign mux_cond_58_shl = {mux_cond_58, 19'h0};
  assign mux_cond_58_pad = mux_cond_58_shl;
  assign mux_cond_59_shl = {mux_cond_59, 2'h0};
  assign mux_cond_59_pad = {17'h0,mux_cond_59_shl};
  assign mux_cond_60_shl = {mux_cond_60, 15'h0};
  assign mux_cond_60_pad = {4'h0,mux_cond_60_shl};
  assign mux_cond_61_shl = {mux_cond_61, 17'h0};
  assign mux_cond_61_pad = {2'h0,mux_cond_61_shl};
  assign mux_cond_62_shl = {mux_cond_62, 11'h0};
  assign mux_cond_62_pad = {8'h0,mux_cond_62_shl};
  assign mux_cond_63_shl = {mux_cond_63, 15'h0};
  assign mux_cond_63_pad = {4'h0,mux_cond_63_shl};
  assign mux_cond_64_shl = {mux_cond_64, 9'h0};
  assign mux_cond_64_pad = {10'h0,mux_cond_64_shl};
  assign mux_cond_65_shl = {mux_cond_65, 17'h0};
  assign mux_cond_65_pad = {2'h0,mux_cond_65_shl};
  assign mux_cond_66_shl = {mux_cond_66, 12'h0};
  assign mux_cond_66_pad = {7'h0,mux_cond_66_shl};
  assign mux_cond_67_shl = {mux_cond_67, 15'h0};
  assign mux_cond_67_pad = {4'h0,mux_cond_67_shl};
  assign mux_cond_68_shl = {mux_cond_68, 17'h0};
  assign mux_cond_68_pad = {2'h0,mux_cond_68_shl};
  assign mux_cond_69_shl = {mux_cond_69, 3'h0};
  assign mux_cond_69_pad = {16'h0,mux_cond_69_shl};
  assign mux_cond_70_shl = {mux_cond_70, 3'h0};
  assign mux_cond_70_pad = {16'h0,mux_cond_70_shl};
  assign sectored_entries_7_valid_1_shl = {sectored_entries_7_valid_1, 12'h0};
  assign sectored_entries_7_valid_1_pad = {7'h0,sectored_entries_7_valid_1_shl};
  assign sectored_entries_5_valid_3_shl = {sectored_entries_5_valid_3, 7'h0};
  assign sectored_entries_5_valid_3_pad = {12'h0,sectored_entries_5_valid_3_shl};
  assign sectored_entries_5_valid_1_shl = {sectored_entries_5_valid_1, 12'h0};
  assign sectored_entries_5_valid_1_pad = {7'h0,sectored_entries_5_valid_1_shl};
  assign sectored_entries_4_valid_1_shl = {sectored_entries_4_valid_1, 12'h0};
  assign sectored_entries_4_valid_1_pad = {7'h0,sectored_entries_4_valid_1_shl};
  assign superpage_entries_0_valid_0_shl = {superpage_entries_0_valid_0, 6'h0};
  assign superpage_entries_0_valid_0_pad = {13'h0,superpage_entries_0_valid_0_shl};
  assign sectored_entries_3_valid_2_shl = {sectored_entries_3_valid_2, 9'h0};
  assign sectored_entries_3_valid_2_pad = {10'h0,sectored_entries_3_valid_2_shl};
  assign sectored_entries_1_valid_0_shl = {sectored_entries_1_valid_0, 9'h0};
  assign sectored_entries_1_valid_0_pad = {10'h0,sectored_entries_1_valid_0_shl};
  assign superpage_entries_3_level_shl = {superpage_entries_3_level, 2'h0};
  assign superpage_entries_3_level_pad = {16'h0,superpage_entries_3_level_shl};
  assign sectored_entries_5_valid_0_shl = {sectored_entries_5_valid_0, 9'h0};
  assign sectored_entries_5_valid_0_pad = {10'h0,sectored_entries_5_valid_0_shl};
  assign sectored_entries_0_valid_1_shl = {sectored_entries_0_valid_1, 12'h0};
  assign sectored_entries_0_valid_1_pad = {7'h0,sectored_entries_0_valid_1_shl};
  assign sectored_entries_3_valid_0_shl = {sectored_entries_3_valid_0, 9'h0};
  assign sectored_entries_3_valid_0_pad = {10'h0,sectored_entries_3_valid_0_shl};
  assign sectored_entries_7_valid_2_shl = {sectored_entries_7_valid_2, 9'h0};
  assign sectored_entries_7_valid_2_pad = {10'h0,sectored_entries_7_valid_2_shl};
  assign sectored_entries_2_valid_3_shl = {sectored_entries_2_valid_3, 7'h0};
  assign sectored_entries_2_valid_3_pad = {12'h0,sectored_entries_2_valid_3_shl};
  assign sectored_entries_4_valid_0_shl = {sectored_entries_4_valid_0, 9'h0};
  assign sectored_entries_4_valid_0_pad = {10'h0,sectored_entries_4_valid_0_shl};
  assign sectored_entries_6_valid_3_shl = {sectored_entries_6_valid_3, 7'h0};
  assign sectored_entries_6_valid_3_pad = {12'h0,sectored_entries_6_valid_3_shl};
  assign sectored_entries_1_valid_3_shl = {sectored_entries_1_valid_3, 7'h0};
  assign sectored_entries_1_valid_3_pad = {12'h0,sectored_entries_1_valid_3_shl};
  assign sectored_entries_6_valid_0_shl = {sectored_entries_6_valid_0, 9'h0};
  assign sectored_entries_6_valid_0_pad = {10'h0,sectored_entries_6_valid_0_shl};
  assign sectored_entries_2_valid_2_shl = {sectored_entries_2_valid_2, 9'h0};
  assign sectored_entries_2_valid_2_pad = {10'h0,sectored_entries_2_valid_2_shl};
  assign sectored_entries_6_valid_2_shl = {sectored_entries_6_valid_2, 9'h0};
  assign sectored_entries_6_valid_2_pad = {10'h0,sectored_entries_6_valid_2_shl};
  assign sectored_entries_6_valid_1_shl = {sectored_entries_6_valid_1, 12'h0};
  assign sectored_entries_6_valid_1_pad = {7'h0,sectored_entries_6_valid_1_shl};
  assign sectored_entries_4_valid_3_shl = {sectored_entries_4_valid_3, 7'h0};
  assign sectored_entries_4_valid_3_pad = {12'h0,sectored_entries_4_valid_3_shl};
  assign sectored_entries_1_valid_2_shl = {sectored_entries_1_valid_2, 9'h0};
  assign sectored_entries_1_valid_2_pad = {10'h0,sectored_entries_1_valid_2_shl};
  assign sectored_entries_5_valid_2_shl = {sectored_entries_5_valid_2, 9'h0};
  assign sectored_entries_5_valid_2_pad = {10'h0,sectored_entries_5_valid_2_shl};
  assign superpage_entries_2_level_shl = {superpage_entries_2_level, 2'h0};
  assign superpage_entries_2_level_pad = {16'h0,superpage_entries_2_level_shl};
  assign superpage_entries_3_valid_0_shl = {superpage_entries_3_valid_0, 6'h0};
  assign superpage_entries_3_valid_0_pad = {13'h0,superpage_entries_3_valid_0_shl};
  assign sectored_entries_1_valid_1_shl = {sectored_entries_1_valid_1, 12'h0};
  assign sectored_entries_1_valid_1_pad = {7'h0,sectored_entries_1_valid_1_shl};
  assign sectored_entries_0_valid_0_shl = {sectored_entries_0_valid_0, 9'h0};
  assign sectored_entries_0_valid_0_pad = {10'h0,sectored_entries_0_valid_0_shl};
  assign superpage_entries_1_valid_0_shl = {superpage_entries_1_valid_0, 6'h0};
  assign superpage_entries_1_valid_0_pad = {13'h0,superpage_entries_1_valid_0_shl};
  assign sectored_entries_0_valid_3_shl = {sectored_entries_0_valid_3, 7'h0};
  assign sectored_entries_0_valid_3_pad = {12'h0,sectored_entries_0_valid_3_shl};
  assign sectored_entries_7_valid_0_shl = {sectored_entries_7_valid_0, 9'h0};
  assign sectored_entries_7_valid_0_pad = {10'h0,sectored_entries_7_valid_0_shl};
  assign sectored_entries_0_valid_2_shl = {sectored_entries_0_valid_2, 9'h0};
  assign sectored_entries_0_valid_2_pad = {10'h0,sectored_entries_0_valid_2_shl};
  assign superpage_entries_0_level_shl = {superpage_entries_0_level, 2'h0};
  assign superpage_entries_0_level_pad = {16'h0,superpage_entries_0_level_shl};
  assign sectored_entries_2_valid_1_shl = {sectored_entries_2_valid_1, 12'h0};
  assign sectored_entries_2_valid_1_pad = {7'h0,sectored_entries_2_valid_1_shl};
  assign sectored_entries_3_valid_1_shl = {sectored_entries_3_valid_1, 12'h0};
  assign sectored_entries_3_valid_1_pad = {7'h0,sectored_entries_3_valid_1_shl};
  assign sectored_entries_2_valid_0_shl = {sectored_entries_2_valid_0, 9'h0};
  assign sectored_entries_2_valid_0_pad = {10'h0,sectored_entries_2_valid_0_shl};
  assign sectored_entries_7_valid_3_shl = {sectored_entries_7_valid_3, 7'h0};
  assign sectored_entries_7_valid_3_pad = {12'h0,sectored_entries_7_valid_3_shl};
  assign sectored_entries_4_valid_2_shl = {sectored_entries_4_valid_2, 9'h0};
  assign sectored_entries_4_valid_2_pad = {10'h0,sectored_entries_4_valid_2_shl};
  assign sectored_entries_3_valid_3_shl = {sectored_entries_3_valid_3, 7'h0};
  assign sectored_entries_3_valid_3_pad = {12'h0,sectored_entries_3_valid_3_shl};
  assign superpage_entries_1_level_shl = {superpage_entries_1_level, 2'h0};
  assign superpage_entries_1_level_pad = {16'h0,superpage_entries_1_level_shl};
  assign superpage_entries_2_valid_0_shl = {superpage_entries_2_valid_0, 6'h0};
  assign superpage_entries_2_valid_0_pad = {13'h0,superpage_entries_2_valid_0_shl};
  assign TLB_1_xor64 = state_pad ^ r_sectored_repl_addr_pad;
  assign TLB_1_xor31 = r_superpage_repl_addr_pad ^ TLB_1_xor64;
  assign TLB_1_xor65 = r_sectored_hit_addr_pad ^ special_entry_valid_0_pad;
  assign TLB_1_xor66 = special_entry_level_pad ^ r_sectored_hit_pad;
  assign TLB_1_xor32 = TLB_1_xor65 ^ TLB_1_xor66;
  assign TLB_1_xor15 = TLB_1_xor31 ^ TLB_1_xor32;
  assign TLB_1_xor68 = mux_cond_1_pad ^ mux_cond_2_pad;
  assign TLB_1_xor33 = mux_cond_0_pad ^ TLB_1_xor68;
  assign TLB_1_xor69 = mux_cond_3_pad ^ mux_cond_4_pad;
  assign TLB_1_xor70 = mux_cond_5_pad ^ mux_cond_6_pad;
  assign TLB_1_xor34 = TLB_1_xor69 ^ TLB_1_xor70;
  assign TLB_1_xor16 = TLB_1_xor33 ^ TLB_1_xor34;
  assign TLB_1_xor7 = TLB_1_xor15 ^ TLB_1_xor16;
  assign TLB_1_xor72 = mux_cond_8_pad ^ mux_cond_9_pad;
  assign TLB_1_xor35 = mux_cond_7_pad ^ TLB_1_xor72;
  assign TLB_1_xor73 = mux_cond_10_pad ^ mux_cond_11_pad;
  assign TLB_1_xor74 = mux_cond_12_pad ^ mux_cond_13_pad;
  assign TLB_1_xor36 = TLB_1_xor73 ^ TLB_1_xor74;
  assign TLB_1_xor17 = TLB_1_xor35 ^ TLB_1_xor36;
  assign TLB_1_xor75 = mux_cond_14_pad ^ mux_cond_15_pad;
  assign TLB_1_xor76 = mux_cond_16_pad ^ mux_cond_17_pad;
  assign TLB_1_xor37 = TLB_1_xor75 ^ TLB_1_xor76;
  assign TLB_1_xor77 = mux_cond_18_pad ^ mux_cond_19_pad;
  assign TLB_1_xor78 = mux_cond_20_pad ^ mux_cond_21_pad;
  assign TLB_1_xor38 = TLB_1_xor77 ^ TLB_1_xor78;
  assign TLB_1_xor18 = TLB_1_xor37 ^ TLB_1_xor38;
  assign TLB_1_xor8 = TLB_1_xor17 ^ TLB_1_xor18;
  assign TLB_1_xor3 = TLB_1_xor7 ^ TLB_1_xor8;
  assign TLB_1_xor80 = mux_cond_23_pad ^ mux_cond_24_pad;
  assign TLB_1_xor39 = mux_cond_22_pad ^ TLB_1_xor80;
  assign TLB_1_xor81 = mux_cond_25_pad ^ mux_cond_26_pad;
  assign TLB_1_xor82 = mux_cond_27_pad ^ mux_cond_28_pad;
  assign TLB_1_xor40 = TLB_1_xor81 ^ TLB_1_xor82;
  assign TLB_1_xor19 = TLB_1_xor39 ^ TLB_1_xor40;
  assign TLB_1_xor83 = mux_cond_29_pad ^ mux_cond_30_pad;
  assign TLB_1_xor84 = mux_cond_31_pad ^ mux_cond_32_pad;
  assign TLB_1_xor41 = TLB_1_xor83 ^ TLB_1_xor84;
  assign TLB_1_xor85 = mux_cond_33_pad ^ mux_cond_34_pad;
  assign TLB_1_xor86 = mux_cond_35_pad ^ mux_cond_36_pad;
  assign TLB_1_xor42 = TLB_1_xor85 ^ TLB_1_xor86;
  assign TLB_1_xor20 = TLB_1_xor41 ^ TLB_1_xor42;
  assign TLB_1_xor9 = TLB_1_xor19 ^ TLB_1_xor20;
  assign TLB_1_xor88 = mux_cond_38_pad ^ mux_cond_39_pad;
  assign TLB_1_xor43 = mux_cond_37_pad ^ TLB_1_xor88;
  assign TLB_1_xor89 = mux_cond_40_pad ^ mux_cond_41_pad;
  assign TLB_1_xor90 = mux_cond_42_pad ^ mux_cond_43_pad;
  assign TLB_1_xor44 = TLB_1_xor89 ^ TLB_1_xor90;
  assign TLB_1_xor21 = TLB_1_xor43 ^ TLB_1_xor44;
  assign TLB_1_xor91 = mux_cond_44_pad ^ mux_cond_45_pad;
  assign TLB_1_xor92 = mux_cond_46_pad ^ mux_cond_47_pad;
  assign TLB_1_xor45 = TLB_1_xor91 ^ TLB_1_xor92;
  assign TLB_1_xor93 = mux_cond_48_pad ^ mux_cond_49_pad;
  assign TLB_1_xor94 = mux_cond_50_pad ^ mux_cond_51_pad;
  assign TLB_1_xor46 = TLB_1_xor93 ^ TLB_1_xor94;
  assign TLB_1_xor22 = TLB_1_xor45 ^ TLB_1_xor46;
  assign TLB_1_xor10 = TLB_1_xor21 ^ TLB_1_xor22;
  assign TLB_1_xor4 = TLB_1_xor9 ^ TLB_1_xor10;
  assign TLB_1_xor1 = TLB_1_xor3 ^ TLB_1_xor4;
  assign TLB_1_xor96 = mux_cond_53_pad ^ mux_cond_54_pad;
  assign TLB_1_xor47 = mux_cond_52_pad ^ TLB_1_xor96;
  assign TLB_1_xor97 = mux_cond_55_pad ^ mux_cond_56_pad;
  assign TLB_1_xor98 = mux_cond_57_pad ^ mux_cond_58_pad;
  assign TLB_1_xor48 = TLB_1_xor97 ^ TLB_1_xor98;
  assign TLB_1_xor23 = TLB_1_xor47 ^ TLB_1_xor48;
  assign TLB_1_xor100 = mux_cond_60_pad ^ mux_cond_61_pad;
  assign TLB_1_xor49 = mux_cond_59_pad ^ TLB_1_xor100;
  assign TLB_1_xor101 = mux_cond_62_pad ^ mux_cond_63_pad;
  assign TLB_1_xor102 = mux_cond_64_pad ^ mux_cond_65_pad;
  assign TLB_1_xor50 = TLB_1_xor101 ^ TLB_1_xor102;
  assign TLB_1_xor24 = TLB_1_xor49 ^ TLB_1_xor50;
  assign TLB_1_xor11 = TLB_1_xor23 ^ TLB_1_xor24;
  assign TLB_1_xor104 = mux_cond_67_pad ^ mux_cond_68_pad;
  assign TLB_1_xor51 = mux_cond_66_pad ^ TLB_1_xor104;
  assign TLB_1_xor105 = mux_cond_69_pad ^ mux_cond_70_pad;
  assign TLB_1_xor106 = sectored_entries_7_valid_1_pad ^ sectored_entries_5_valid_3_pad;
  assign TLB_1_xor52 = TLB_1_xor105 ^ TLB_1_xor106;
  assign TLB_1_xor25 = TLB_1_xor51 ^ TLB_1_xor52;
  assign TLB_1_xor107 = sectored_entries_5_valid_1_pad ^ sectored_entries_4_valid_1_pad;
  assign TLB_1_xor108 = superpage_entries_0_valid_0_pad ^ sectored_entries_3_valid_2_pad;
  assign TLB_1_xor53 = TLB_1_xor107 ^ TLB_1_xor108;
  assign TLB_1_xor109 = sectored_entries_1_valid_0_pad ^ superpage_entries_3_level_pad;
  assign TLB_1_xor110 = sectored_entries_5_valid_0_pad ^ sectored_entries_0_valid_1_pad;
  assign TLB_1_xor54 = TLB_1_xor109 ^ TLB_1_xor110;
  assign TLB_1_xor26 = TLB_1_xor53 ^ TLB_1_xor54;
  assign TLB_1_xor12 = TLB_1_xor25 ^ TLB_1_xor26;
  assign TLB_1_xor5 = TLB_1_xor11 ^ TLB_1_xor12;
  assign TLB_1_xor112 = sectored_entries_7_valid_2_pad ^ sectored_entries_2_valid_3_pad;
  assign TLB_1_xor55 = sectored_entries_3_valid_0_pad ^ TLB_1_xor112;
  assign TLB_1_xor113 = sectored_entries_4_valid_0_pad ^ sectored_entries_6_valid_3_pad;
  assign TLB_1_xor114 = sectored_entries_1_valid_3_pad ^ sectored_entries_6_valid_0_pad;
  assign TLB_1_xor56 = TLB_1_xor113 ^ TLB_1_xor114;
  assign TLB_1_xor27 = TLB_1_xor55 ^ TLB_1_xor56;
  assign TLB_1_xor115 = sectored_entries_2_valid_2_pad ^ sectored_entries_6_valid_2_pad;
  assign TLB_1_xor116 = sectored_entries_6_valid_1_pad ^ sectored_entries_4_valid_3_pad;
  assign TLB_1_xor57 = TLB_1_xor115 ^ TLB_1_xor116;
  assign TLB_1_xor117 = sectored_entries_1_valid_2_pad ^ sectored_entries_5_valid_2_pad;
  assign TLB_1_xor118 = superpage_entries_2_level_pad ^ superpage_entries_3_valid_0_pad;
  assign TLB_1_xor58 = TLB_1_xor117 ^ TLB_1_xor118;
  assign TLB_1_xor28 = TLB_1_xor57 ^ TLB_1_xor58;
  assign TLB_1_xor13 = TLB_1_xor27 ^ TLB_1_xor28;
  assign TLB_1_xor120 = sectored_entries_0_valid_0_pad ^ superpage_entries_1_valid_0_pad;
  assign TLB_1_xor59 = sectored_entries_1_valid_1_pad ^ TLB_1_xor120;
  assign TLB_1_xor121 = sectored_entries_0_valid_3_pad ^ sectored_entries_7_valid_0_pad;
  assign TLB_1_xor122 = sectored_entries_0_valid_2_pad ^ superpage_entries_0_level_pad;
  assign TLB_1_xor60 = TLB_1_xor121 ^ TLB_1_xor122;
  assign TLB_1_xor29 = TLB_1_xor59 ^ TLB_1_xor60;
  assign TLB_1_xor123 = sectored_entries_2_valid_1_pad ^ sectored_entries_3_valid_1_pad;
  assign TLB_1_xor124 = sectored_entries_2_valid_0_pad ^ sectored_entries_7_valid_3_pad;
  assign TLB_1_xor61 = TLB_1_xor123 ^ TLB_1_xor124;
  assign TLB_1_xor125 = sectored_entries_4_valid_2_pad ^ sectored_entries_3_valid_3_pad;
  assign TLB_1_xor126 = superpage_entries_1_level_pad ^ superpage_entries_2_valid_0_pad;
  assign TLB_1_xor62 = TLB_1_xor125 ^ TLB_1_xor126;
  assign TLB_1_xor30 = TLB_1_xor61 ^ TLB_1_xor62;
  assign TLB_1_xor14 = TLB_1_xor29 ^ TLB_1_xor30;
  assign TLB_1_xor6 = TLB_1_xor13 ^ TLB_1_xor14;
  assign TLB_1_xor2 = TLB_1_xor5 ^ TLB_1_xor6;
  assign TLB_1_xor0 = TLB_1_xor1 ^ TLB_1_xor2;
  assign pmp_sum = TLB_1_covSum + pmp_io_covSum;
  assign io_covSum = pmp_sum;
  assign stopEn0 = io_sfence_valid & ~_T_2949;
  assign pmp_metaAssert_wire = pmp_metaAssert;
  assign TLB_1_or0 = stopEn0 | pmp_metaAssert_wire;
  assign metaAssert = TLB_1_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sectored_entries_0_tag = _RAND_0[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  sectored_entries_0_data_0 = _RAND_1[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  sectored_entries_0_data_1 = _RAND_2[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{`RANDOM}};
  sectored_entries_0_data_2 = _RAND_3[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{`RANDOM}};
  sectored_entries_0_data_3 = _RAND_4[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  sectored_entries_0_valid_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sectored_entries_0_valid_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  sectored_entries_0_valid_2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sectored_entries_0_valid_3 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  sectored_entries_1_tag = _RAND_9[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {2{`RANDOM}};
  sectored_entries_1_data_0 = _RAND_10[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{`RANDOM}};
  sectored_entries_1_data_1 = _RAND_11[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {2{`RANDOM}};
  sectored_entries_1_data_2 = _RAND_12[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  sectored_entries_1_data_3 = _RAND_13[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  sectored_entries_1_valid_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  sectored_entries_1_valid_1 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  sectored_entries_1_valid_2 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  sectored_entries_1_valid_3 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  sectored_entries_2_tag = _RAND_18[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{`RANDOM}};
  sectored_entries_2_data_0 = _RAND_19[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{`RANDOM}};
  sectored_entries_2_data_1 = _RAND_20[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{`RANDOM}};
  sectored_entries_2_data_2 = _RAND_21[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {2{`RANDOM}};
  sectored_entries_2_data_3 = _RAND_22[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  sectored_entries_2_valid_0 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  sectored_entries_2_valid_1 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  sectored_entries_2_valid_2 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  sectored_entries_2_valid_3 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  sectored_entries_3_tag = _RAND_27[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {2{`RANDOM}};
  sectored_entries_3_data_0 = _RAND_28[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {2{`RANDOM}};
  sectored_entries_3_data_1 = _RAND_29[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {2{`RANDOM}};
  sectored_entries_3_data_2 = _RAND_30[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{`RANDOM}};
  sectored_entries_3_data_3 = _RAND_31[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  sectored_entries_3_valid_0 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  sectored_entries_3_valid_1 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  sectored_entries_3_valid_2 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  sectored_entries_3_valid_3 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  sectored_entries_4_tag = _RAND_36[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{`RANDOM}};
  sectored_entries_4_data_0 = _RAND_37[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {2{`RANDOM}};
  sectored_entries_4_data_1 = _RAND_38[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{`RANDOM}};
  sectored_entries_4_data_2 = _RAND_39[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {2{`RANDOM}};
  sectored_entries_4_data_3 = _RAND_40[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  sectored_entries_4_valid_0 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  sectored_entries_4_valid_1 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  sectored_entries_4_valid_2 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  sectored_entries_4_valid_3 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  sectored_entries_5_tag = _RAND_45[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {2{`RANDOM}};
  sectored_entries_5_data_0 = _RAND_46[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {2{`RANDOM}};
  sectored_entries_5_data_1 = _RAND_47[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {2{`RANDOM}};
  sectored_entries_5_data_2 = _RAND_48[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {2{`RANDOM}};
  sectored_entries_5_data_3 = _RAND_49[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  sectored_entries_5_valid_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  sectored_entries_5_valid_1 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  sectored_entries_5_valid_2 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  sectored_entries_5_valid_3 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  sectored_entries_6_tag = _RAND_54[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {2{`RANDOM}};
  sectored_entries_6_data_0 = _RAND_55[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {2{`RANDOM}};
  sectored_entries_6_data_1 = _RAND_56[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {2{`RANDOM}};
  sectored_entries_6_data_2 = _RAND_57[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {2{`RANDOM}};
  sectored_entries_6_data_3 = _RAND_58[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  sectored_entries_6_valid_0 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  sectored_entries_6_valid_1 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  sectored_entries_6_valid_2 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  sectored_entries_6_valid_3 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  sectored_entries_7_tag = _RAND_63[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {2{`RANDOM}};
  sectored_entries_7_data_0 = _RAND_64[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {2{`RANDOM}};
  sectored_entries_7_data_1 = _RAND_65[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {2{`RANDOM}};
  sectored_entries_7_data_2 = _RAND_66[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {2{`RANDOM}};
  sectored_entries_7_data_3 = _RAND_67[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  sectored_entries_7_valid_0 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  sectored_entries_7_valid_1 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  sectored_entries_7_valid_2 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  sectored_entries_7_valid_3 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  superpage_entries_0_level = _RAND_72[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  superpage_entries_0_tag = _RAND_73[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {2{`RANDOM}};
  superpage_entries_0_data_0 = _RAND_74[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  superpage_entries_0_valid_0 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  superpage_entries_1_level = _RAND_76[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  superpage_entries_1_tag = _RAND_77[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {2{`RANDOM}};
  superpage_entries_1_data_0 = _RAND_78[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  superpage_entries_1_valid_0 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  superpage_entries_2_level = _RAND_80[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  superpage_entries_2_tag = _RAND_81[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {2{`RANDOM}};
  superpage_entries_2_data_0 = _RAND_82[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  superpage_entries_2_valid_0 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  superpage_entries_3_level = _RAND_84[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  superpage_entries_3_tag = _RAND_85[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {2{`RANDOM}};
  superpage_entries_3_data_0 = _RAND_86[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  superpage_entries_3_valid_0 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  special_entry_level = _RAND_88[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  special_entry_tag = _RAND_89[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {2{`RANDOM}};
  special_entry_data_0 = _RAND_90[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  special_entry_valid_0 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  state = _RAND_92[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  r_refill_tag = _RAND_93[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  r_superpage_repl_addr = _RAND_94[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  r_sectored_repl_addr = _RAND_95[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  r_sectored_hit_addr = _RAND_96[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  r_sectored_hit = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  vpoffset_cfg_value = _RAND_98[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  requestedVPN = _RAND_99[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_2554 = _RAND_100[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_2556 = _RAND_101[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  TLB_1_state = _RAND_102[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    TLB_1_cov[initvar] = _RAND_103[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  TLB_1_covSum = _RAND_104[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  TLB_1_metaAssert = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      sectored_entries_0_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1505) begin
            sectored_entries_0_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1505) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_0 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_data_1 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1505) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_1 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_data_2 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1505) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_2 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_data_3 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1505) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_3 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_0_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2957) begin
          if (sectored_entries_0_data_0[0]) begin
            sectored_entries_0_valid_0 <= 1'h0;
          end else if (_T_727) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_0_valid_0 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1505) begin
                    sectored_entries_0_valid_0 <= _GEN_85;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1505) begin
                  sectored_entries_0_valid_0 <= _GEN_85;
                end
              end
            end
          end
        end else if (_T_727) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_0_valid_0 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1505) begin
                  sectored_entries_0_valid_0 <= _GEN_85;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1505) begin
                sectored_entries_0_valid_0 <= _GEN_85;
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_0 <= _GEN_656;
      end
    end else begin
      sectored_entries_0_valid_0 <= _GEN_473;
    end
    if (metaReset) begin
      sectored_entries_0_valid_1 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_0_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2957) begin
          if (sectored_entries_0_data_1[0]) begin
            sectored_entries_0_valid_1 <= 1'h0;
          end else if (_T_727) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_0_valid_1 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1505) begin
                    sectored_entries_0_valid_1 <= _GEN_86;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1505) begin
                  sectored_entries_0_valid_1 <= _GEN_86;
                end
              end
            end
          end
        end else if (_T_727) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_0_valid_1 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1505) begin
                  sectored_entries_0_valid_1 <= _GEN_86;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1505) begin
                sectored_entries_0_valid_1 <= _GEN_86;
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_1 <= _GEN_657;
      end
    end else begin
      sectored_entries_0_valid_1 <= _GEN_474;
    end
    if (metaReset) begin
      sectored_entries_0_valid_2 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_0_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2957) begin
          if (sectored_entries_0_data_2[0]) begin
            sectored_entries_0_valid_2 <= 1'h0;
          end else if (_T_727) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_0_valid_2 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1505) begin
                    sectored_entries_0_valid_2 <= _GEN_87;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1505) begin
                  sectored_entries_0_valid_2 <= _GEN_87;
                end
              end
            end
          end
        end else if (_T_727) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_0_valid_2 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1505) begin
                  sectored_entries_0_valid_2 <= _GEN_87;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1505) begin
                sectored_entries_0_valid_2 <= _GEN_87;
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_2 <= _GEN_658;
      end
    end else begin
      sectored_entries_0_valid_2 <= _GEN_475;
    end
    if (metaReset) begin
      sectored_entries_0_valid_3 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_0_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2957) begin
          if (sectored_entries_0_data_3[0]) begin
            sectored_entries_0_valid_3 <= 1'h0;
          end else if (_T_727) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_0_valid_3 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1505) begin
                    sectored_entries_0_valid_3 <= _GEN_88;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1505) begin
                  sectored_entries_0_valid_3 <= _GEN_88;
                end
              end
            end
          end
        end else if (_T_727) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_0_valid_3 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1505) begin
                  sectored_entries_0_valid_3 <= _GEN_88;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1505) begin
                sectored_entries_0_valid_3 <= _GEN_88;
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_3 <= _GEN_659;
      end
    end else begin
      sectored_entries_0_valid_3 <= _GEN_476;
    end
    if (metaReset) begin
      sectored_entries_1_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1522) begin
            sectored_entries_1_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_1_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1522) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_0 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_1_data_1 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1522) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_1 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_1_data_2 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1522) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_2 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_1_data_3 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1522) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_3 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_1_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_1_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3128) begin
          if (sectored_entries_1_data_0[0]) begin
            sectored_entries_1_valid_0 <= 1'h0;
          end else if (_T_733) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_1_valid_0 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1522) begin
                    sectored_entries_1_valid_0 <= _GEN_107;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1522) begin
                  sectored_entries_1_valid_0 <= _GEN_107;
                end
              end
            end
          end
        end else if (_T_733) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_1_valid_0 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1522) begin
                  sectored_entries_1_valid_0 <= _GEN_107;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1522) begin
                sectored_entries_1_valid_0 <= _GEN_107;
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_0 <= _GEN_684;
      end
    end else begin
      sectored_entries_1_valid_0 <= _GEN_483;
    end
    if (metaReset) begin
      sectored_entries_1_valid_1 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_1_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3128) begin
          if (sectored_entries_1_data_1[0]) begin
            sectored_entries_1_valid_1 <= 1'h0;
          end else if (_T_733) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_1_valid_1 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1522) begin
                    sectored_entries_1_valid_1 <= _GEN_108;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1522) begin
                  sectored_entries_1_valid_1 <= _GEN_108;
                end
              end
            end
          end
        end else if (_T_733) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_1_valid_1 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1522) begin
                  sectored_entries_1_valid_1 <= _GEN_108;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1522) begin
                sectored_entries_1_valid_1 <= _GEN_108;
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_1 <= _GEN_685;
      end
    end else begin
      sectored_entries_1_valid_1 <= _GEN_484;
    end
    if (metaReset) begin
      sectored_entries_1_valid_2 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_1_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3128) begin
          if (sectored_entries_1_data_2[0]) begin
            sectored_entries_1_valid_2 <= 1'h0;
          end else if (_T_733) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_1_valid_2 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1522) begin
                    sectored_entries_1_valid_2 <= _GEN_109;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1522) begin
                  sectored_entries_1_valid_2 <= _GEN_109;
                end
              end
            end
          end
        end else if (_T_733) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_1_valid_2 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1522) begin
                  sectored_entries_1_valid_2 <= _GEN_109;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1522) begin
                sectored_entries_1_valid_2 <= _GEN_109;
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_2 <= _GEN_686;
      end
    end else begin
      sectored_entries_1_valid_2 <= _GEN_485;
    end
    if (metaReset) begin
      sectored_entries_1_valid_3 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_1_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3128) begin
          if (sectored_entries_1_data_3[0]) begin
            sectored_entries_1_valid_3 <= 1'h0;
          end else if (_T_733) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_1_valid_3 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1522) begin
                    sectored_entries_1_valid_3 <= _GEN_110;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1522) begin
                  sectored_entries_1_valid_3 <= _GEN_110;
                end
              end
            end
          end
        end else if (_T_733) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_1_valid_3 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1522) begin
                  sectored_entries_1_valid_3 <= _GEN_110;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1522) begin
                sectored_entries_1_valid_3 <= _GEN_110;
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_3 <= _GEN_687;
      end
    end else begin
      sectored_entries_1_valid_3 <= _GEN_486;
    end
    if (metaReset) begin
      sectored_entries_2_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1539) begin
            sectored_entries_2_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_2_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1539) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_0 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_2_data_1 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1539) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_1 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_2_data_2 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1539) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_2 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_2_data_3 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1539) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_3 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_2_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_2_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3299) begin
          if (sectored_entries_2_data_0[0]) begin
            sectored_entries_2_valid_0 <= 1'h0;
          end else if (_T_739) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_2_valid_0 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1539) begin
                    sectored_entries_2_valid_0 <= _GEN_129;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1539) begin
                  sectored_entries_2_valid_0 <= _GEN_129;
                end
              end
            end
          end
        end else if (_T_739) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_2_valid_0 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1539) begin
                  sectored_entries_2_valid_0 <= _GEN_129;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1539) begin
                sectored_entries_2_valid_0 <= _GEN_129;
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_0 <= _GEN_712;
      end
    end else begin
      sectored_entries_2_valid_0 <= _GEN_493;
    end
    if (metaReset) begin
      sectored_entries_2_valid_1 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_2_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3299) begin
          if (sectored_entries_2_data_1[0]) begin
            sectored_entries_2_valid_1 <= 1'h0;
          end else if (_T_739) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_2_valid_1 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1539) begin
                    sectored_entries_2_valid_1 <= _GEN_130;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1539) begin
                  sectored_entries_2_valid_1 <= _GEN_130;
                end
              end
            end
          end
        end else if (_T_739) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_2_valid_1 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1539) begin
                  sectored_entries_2_valid_1 <= _GEN_130;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1539) begin
                sectored_entries_2_valid_1 <= _GEN_130;
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_1 <= _GEN_713;
      end
    end else begin
      sectored_entries_2_valid_1 <= _GEN_494;
    end
    if (metaReset) begin
      sectored_entries_2_valid_2 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_2_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3299) begin
          if (sectored_entries_2_data_2[0]) begin
            sectored_entries_2_valid_2 <= 1'h0;
          end else if (_T_739) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_2_valid_2 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1539) begin
                    sectored_entries_2_valid_2 <= _GEN_131;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1539) begin
                  sectored_entries_2_valid_2 <= _GEN_131;
                end
              end
            end
          end
        end else if (_T_739) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_2_valid_2 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1539) begin
                  sectored_entries_2_valid_2 <= _GEN_131;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1539) begin
                sectored_entries_2_valid_2 <= _GEN_131;
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_2 <= _GEN_714;
      end
    end else begin
      sectored_entries_2_valid_2 <= _GEN_495;
    end
    if (metaReset) begin
      sectored_entries_2_valid_3 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_2_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3299) begin
          if (sectored_entries_2_data_3[0]) begin
            sectored_entries_2_valid_3 <= 1'h0;
          end else if (_T_739) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_2_valid_3 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1539) begin
                    sectored_entries_2_valid_3 <= _GEN_132;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1539) begin
                  sectored_entries_2_valid_3 <= _GEN_132;
                end
              end
            end
          end
        end else if (_T_739) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_2_valid_3 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1539) begin
                  sectored_entries_2_valid_3 <= _GEN_132;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1539) begin
                sectored_entries_2_valid_3 <= _GEN_132;
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_3 <= _GEN_715;
      end
    end else begin
      sectored_entries_2_valid_3 <= _GEN_496;
    end
    if (metaReset) begin
      sectored_entries_3_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1556) begin
            sectored_entries_3_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_3_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1556) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_0 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_3_data_1 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1556) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_1 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_3_data_2 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1556) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_2 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_3_data_3 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1556) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_3 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_3_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_3_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3470) begin
          if (sectored_entries_3_data_0[0]) begin
            sectored_entries_3_valid_0 <= 1'h0;
          end else if (_T_745) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_3_valid_0 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1556) begin
                    sectored_entries_3_valid_0 <= _GEN_151;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1556) begin
                  sectored_entries_3_valid_0 <= _GEN_151;
                end
              end
            end
          end
        end else if (_T_745) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_3_valid_0 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1556) begin
                  sectored_entries_3_valid_0 <= _GEN_151;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1556) begin
                sectored_entries_3_valid_0 <= _GEN_151;
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_0 <= _GEN_740;
      end
    end else begin
      sectored_entries_3_valid_0 <= _GEN_503;
    end
    if (metaReset) begin
      sectored_entries_3_valid_1 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_3_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3470) begin
          if (sectored_entries_3_data_1[0]) begin
            sectored_entries_3_valid_1 <= 1'h0;
          end else if (_T_745) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_3_valid_1 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1556) begin
                    sectored_entries_3_valid_1 <= _GEN_152;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1556) begin
                  sectored_entries_3_valid_1 <= _GEN_152;
                end
              end
            end
          end
        end else if (_T_745) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_3_valid_1 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1556) begin
                  sectored_entries_3_valid_1 <= _GEN_152;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1556) begin
                sectored_entries_3_valid_1 <= _GEN_152;
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_1 <= _GEN_741;
      end
    end else begin
      sectored_entries_3_valid_1 <= _GEN_504;
    end
    if (metaReset) begin
      sectored_entries_3_valid_2 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_3_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3470) begin
          if (sectored_entries_3_data_2[0]) begin
            sectored_entries_3_valid_2 <= 1'h0;
          end else if (_T_745) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_3_valid_2 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1556) begin
                    sectored_entries_3_valid_2 <= _GEN_153;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1556) begin
                  sectored_entries_3_valid_2 <= _GEN_153;
                end
              end
            end
          end
        end else if (_T_745) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_3_valid_2 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1556) begin
                  sectored_entries_3_valid_2 <= _GEN_153;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1556) begin
                sectored_entries_3_valid_2 <= _GEN_153;
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_2 <= _GEN_742;
      end
    end else begin
      sectored_entries_3_valid_2 <= _GEN_505;
    end
    if (metaReset) begin
      sectored_entries_3_valid_3 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_3_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3470) begin
          if (sectored_entries_3_data_3[0]) begin
            sectored_entries_3_valid_3 <= 1'h0;
          end else if (_T_745) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_3_valid_3 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1556) begin
                    sectored_entries_3_valid_3 <= _GEN_154;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1556) begin
                  sectored_entries_3_valid_3 <= _GEN_154;
                end
              end
            end
          end
        end else if (_T_745) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_3_valid_3 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1556) begin
                  sectored_entries_3_valid_3 <= _GEN_154;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1556) begin
                sectored_entries_3_valid_3 <= _GEN_154;
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_3 <= _GEN_743;
      end
    end else begin
      sectored_entries_3_valid_3 <= _GEN_506;
    end
    if (metaReset) begin
      sectored_entries_4_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1573) begin
            sectored_entries_4_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_4_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1573) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_0 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_4_data_1 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1573) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_1 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_4_data_2 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1573) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_2 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_4_data_3 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1573) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_3 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_4_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_4_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3641) begin
          if (sectored_entries_4_data_0[0]) begin
            sectored_entries_4_valid_0 <= 1'h0;
          end else if (_T_751) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_4_valid_0 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1573) begin
                    sectored_entries_4_valid_0 <= _GEN_173;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1573) begin
                  sectored_entries_4_valid_0 <= _GEN_173;
                end
              end
            end
          end
        end else if (_T_751) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_4_valid_0 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1573) begin
                  sectored_entries_4_valid_0 <= _GEN_173;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1573) begin
                sectored_entries_4_valid_0 <= _GEN_173;
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_0 <= _GEN_768;
      end
    end else begin
      sectored_entries_4_valid_0 <= _GEN_513;
    end
    if (metaReset) begin
      sectored_entries_4_valid_1 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_4_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3641) begin
          if (sectored_entries_4_data_1[0]) begin
            sectored_entries_4_valid_1 <= 1'h0;
          end else if (_T_751) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_4_valid_1 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1573) begin
                    sectored_entries_4_valid_1 <= _GEN_174;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1573) begin
                  sectored_entries_4_valid_1 <= _GEN_174;
                end
              end
            end
          end
        end else if (_T_751) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_4_valid_1 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1573) begin
                  sectored_entries_4_valid_1 <= _GEN_174;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1573) begin
                sectored_entries_4_valid_1 <= _GEN_174;
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_1 <= _GEN_769;
      end
    end else begin
      sectored_entries_4_valid_1 <= _GEN_514;
    end
    if (metaReset) begin
      sectored_entries_4_valid_2 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_4_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3641) begin
          if (sectored_entries_4_data_2[0]) begin
            sectored_entries_4_valid_2 <= 1'h0;
          end else if (_T_751) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_4_valid_2 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1573) begin
                    sectored_entries_4_valid_2 <= _GEN_175;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1573) begin
                  sectored_entries_4_valid_2 <= _GEN_175;
                end
              end
            end
          end
        end else if (_T_751) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_4_valid_2 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1573) begin
                  sectored_entries_4_valid_2 <= _GEN_175;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1573) begin
                sectored_entries_4_valid_2 <= _GEN_175;
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_2 <= _GEN_770;
      end
    end else begin
      sectored_entries_4_valid_2 <= _GEN_515;
    end
    if (metaReset) begin
      sectored_entries_4_valid_3 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_4_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3641) begin
          if (sectored_entries_4_data_3[0]) begin
            sectored_entries_4_valid_3 <= 1'h0;
          end else if (_T_751) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_4_valid_3 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1573) begin
                    sectored_entries_4_valid_3 <= _GEN_176;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1573) begin
                  sectored_entries_4_valid_3 <= _GEN_176;
                end
              end
            end
          end
        end else if (_T_751) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_4_valid_3 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1573) begin
                  sectored_entries_4_valid_3 <= _GEN_176;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1573) begin
                sectored_entries_4_valid_3 <= _GEN_176;
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_3 <= _GEN_771;
      end
    end else begin
      sectored_entries_4_valid_3 <= _GEN_516;
    end
    if (metaReset) begin
      sectored_entries_5_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1590) begin
            sectored_entries_5_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_5_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1590) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_0 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_5_data_1 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1590) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_1 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_5_data_2 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1590) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_2 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_5_data_3 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1590) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_3 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_5_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_5_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3812) begin
          if (sectored_entries_5_data_0[0]) begin
            sectored_entries_5_valid_0 <= 1'h0;
          end else if (_T_757) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_5_valid_0 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1590) begin
                    sectored_entries_5_valid_0 <= _GEN_195;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1590) begin
                  sectored_entries_5_valid_0 <= _GEN_195;
                end
              end
            end
          end
        end else if (_T_757) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_5_valid_0 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1590) begin
                  sectored_entries_5_valid_0 <= _GEN_195;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1590) begin
                sectored_entries_5_valid_0 <= _GEN_195;
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_0 <= _GEN_796;
      end
    end else begin
      sectored_entries_5_valid_0 <= _GEN_523;
    end
    if (metaReset) begin
      sectored_entries_5_valid_1 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_5_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3812) begin
          if (sectored_entries_5_data_1[0]) begin
            sectored_entries_5_valid_1 <= 1'h0;
          end else if (_T_757) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_5_valid_1 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1590) begin
                    sectored_entries_5_valid_1 <= _GEN_196;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1590) begin
                  sectored_entries_5_valid_1 <= _GEN_196;
                end
              end
            end
          end
        end else if (_T_757) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_5_valid_1 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1590) begin
                  sectored_entries_5_valid_1 <= _GEN_196;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1590) begin
                sectored_entries_5_valid_1 <= _GEN_196;
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_1 <= _GEN_797;
      end
    end else begin
      sectored_entries_5_valid_1 <= _GEN_524;
    end
    if (metaReset) begin
      sectored_entries_5_valid_2 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_5_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3812) begin
          if (sectored_entries_5_data_2[0]) begin
            sectored_entries_5_valid_2 <= 1'h0;
          end else if (_T_757) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_5_valid_2 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1590) begin
                    sectored_entries_5_valid_2 <= _GEN_197;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1590) begin
                  sectored_entries_5_valid_2 <= _GEN_197;
                end
              end
            end
          end
        end else if (_T_757) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_5_valid_2 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1590) begin
                  sectored_entries_5_valid_2 <= _GEN_197;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1590) begin
                sectored_entries_5_valid_2 <= _GEN_197;
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_2 <= _GEN_798;
      end
    end else begin
      sectored_entries_5_valid_2 <= _GEN_525;
    end
    if (metaReset) begin
      sectored_entries_5_valid_3 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_5_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3812) begin
          if (sectored_entries_5_data_3[0]) begin
            sectored_entries_5_valid_3 <= 1'h0;
          end else if (_T_757) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_5_valid_3 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1590) begin
                    sectored_entries_5_valid_3 <= _GEN_198;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1590) begin
                  sectored_entries_5_valid_3 <= _GEN_198;
                end
              end
            end
          end
        end else if (_T_757) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_5_valid_3 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1590) begin
                  sectored_entries_5_valid_3 <= _GEN_198;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1590) begin
                sectored_entries_5_valid_3 <= _GEN_198;
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_3 <= _GEN_799;
      end
    end else begin
      sectored_entries_5_valid_3 <= _GEN_526;
    end
    if (metaReset) begin
      sectored_entries_6_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1607) begin
            sectored_entries_6_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_6_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1607) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_0 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_6_data_1 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1607) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_1 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_6_data_2 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1607) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_2 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_6_data_3 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1607) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_3 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_6_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_6_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3983) begin
          if (sectored_entries_6_data_0[0]) begin
            sectored_entries_6_valid_0 <= 1'h0;
          end else if (_T_763) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_6_valid_0 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1607) begin
                    sectored_entries_6_valid_0 <= _GEN_217;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1607) begin
                  sectored_entries_6_valid_0 <= _GEN_217;
                end
              end
            end
          end
        end else if (_T_763) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_6_valid_0 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1607) begin
                  sectored_entries_6_valid_0 <= _GEN_217;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1607) begin
                sectored_entries_6_valid_0 <= _GEN_217;
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_0 <= _GEN_824;
      end
    end else begin
      sectored_entries_6_valid_0 <= _GEN_533;
    end
    if (metaReset) begin
      sectored_entries_6_valid_1 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_6_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3983) begin
          if (sectored_entries_6_data_1[0]) begin
            sectored_entries_6_valid_1 <= 1'h0;
          end else if (_T_763) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_6_valid_1 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1607) begin
                    sectored_entries_6_valid_1 <= _GEN_218;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1607) begin
                  sectored_entries_6_valid_1 <= _GEN_218;
                end
              end
            end
          end
        end else if (_T_763) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_6_valid_1 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1607) begin
                  sectored_entries_6_valid_1 <= _GEN_218;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1607) begin
                sectored_entries_6_valid_1 <= _GEN_218;
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_1 <= _GEN_825;
      end
    end else begin
      sectored_entries_6_valid_1 <= _GEN_534;
    end
    if (metaReset) begin
      sectored_entries_6_valid_2 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_6_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3983) begin
          if (sectored_entries_6_data_2[0]) begin
            sectored_entries_6_valid_2 <= 1'h0;
          end else if (_T_763) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_6_valid_2 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1607) begin
                    sectored_entries_6_valid_2 <= _GEN_219;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1607) begin
                  sectored_entries_6_valid_2 <= _GEN_219;
                end
              end
            end
          end
        end else if (_T_763) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_6_valid_2 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1607) begin
                  sectored_entries_6_valid_2 <= _GEN_219;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1607) begin
                sectored_entries_6_valid_2 <= _GEN_219;
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_2 <= _GEN_826;
      end
    end else begin
      sectored_entries_6_valid_2 <= _GEN_535;
    end
    if (metaReset) begin
      sectored_entries_6_valid_3 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_6_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3983) begin
          if (sectored_entries_6_data_3[0]) begin
            sectored_entries_6_valid_3 <= 1'h0;
          end else if (_T_763) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_6_valid_3 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1607) begin
                    sectored_entries_6_valid_3 <= _GEN_220;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1607) begin
                  sectored_entries_6_valid_3 <= _GEN_220;
                end
              end
            end
          end
        end else if (_T_763) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_6_valid_3 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1607) begin
                  sectored_entries_6_valid_3 <= _GEN_220;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1607) begin
                sectored_entries_6_valid_3 <= _GEN_220;
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_3 <= _GEN_827;
      end
    end else begin
      sectored_entries_6_valid_3 <= _GEN_536;
    end
    if (metaReset) begin
      sectored_entries_7_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1624) begin
            sectored_entries_7_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_7_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1624) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_0 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_7_data_1 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1624) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_1 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_7_data_2 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1624) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_2 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_7_data_3 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_1439)) begin
          if (_T_1624) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_3 <= _T_1438;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_7_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_7_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_4154) begin
          if (sectored_entries_7_data_0[0]) begin
            sectored_entries_7_valid_0 <= 1'h0;
          end else if (_T_769) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_7_valid_0 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1624) begin
                    sectored_entries_7_valid_0 <= _GEN_239;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1624) begin
                  sectored_entries_7_valid_0 <= _GEN_239;
                end
              end
            end
          end
        end else if (_T_769) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_7_valid_0 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1624) begin
                  sectored_entries_7_valid_0 <= _GEN_239;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1624) begin
                sectored_entries_7_valid_0 <= _GEN_239;
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_0 <= _GEN_852;
      end
    end else begin
      sectored_entries_7_valid_0 <= _GEN_543;
    end
    if (metaReset) begin
      sectored_entries_7_valid_1 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_7_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_4154) begin
          if (sectored_entries_7_data_1[0]) begin
            sectored_entries_7_valid_1 <= 1'h0;
          end else if (_T_769) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_7_valid_1 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1624) begin
                    sectored_entries_7_valid_1 <= _GEN_240;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1624) begin
                  sectored_entries_7_valid_1 <= _GEN_240;
                end
              end
            end
          end
        end else if (_T_769) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_7_valid_1 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1624) begin
                  sectored_entries_7_valid_1 <= _GEN_240;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1624) begin
                sectored_entries_7_valid_1 <= _GEN_240;
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_1 <= _GEN_853;
      end
    end else begin
      sectored_entries_7_valid_1 <= _GEN_544;
    end
    if (metaReset) begin
      sectored_entries_7_valid_2 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_7_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_4154) begin
          if (sectored_entries_7_data_2[0]) begin
            sectored_entries_7_valid_2 <= 1'h0;
          end else if (_T_769) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_7_valid_2 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1624) begin
                    sectored_entries_7_valid_2 <= _GEN_241;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1624) begin
                  sectored_entries_7_valid_2 <= _GEN_241;
                end
              end
            end
          end
        end else if (_T_769) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_7_valid_2 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1624) begin
                  sectored_entries_7_valid_2 <= _GEN_241;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1624) begin
                sectored_entries_7_valid_2 <= _GEN_241;
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_2 <= _GEN_854;
      end
    end else begin
      sectored_entries_7_valid_2 <= _GEN_545;
    end
    if (metaReset) begin
      sectored_entries_7_valid_3 <= 1'h0;
    end else if (_T_4530) begin
      sectored_entries_7_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_4154) begin
          if (sectored_entries_7_data_3[0]) begin
            sectored_entries_7_valid_3 <= 1'h0;
          end else if (_T_769) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_7_valid_3 <= 1'h0;
            end else if (_T_1385) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_1439)) begin
                  if (_T_1624) begin
                    sectored_entries_7_valid_3 <= _GEN_242;
                  end
                end
              end
            end
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1624) begin
                  sectored_entries_7_valid_3 <= _GEN_242;
                end
              end
            end
          end
        end else if (_T_769) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_7_valid_3 <= 1'h0;
          end else if (_T_1385) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_1439)) begin
                if (_T_1624) begin
                  sectored_entries_7_valid_3 <= _GEN_242;
                end
              end
            end
          end
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_1439)) begin
              if (_T_1624) begin
                sectored_entries_7_valid_3 <= _GEN_242;
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_3 <= _GEN_855;
      end
    end else begin
      sectored_entries_7_valid_3 <= _GEN_546;
    end
    if (metaReset) begin
      superpage_entries_0_level <= 2'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1440) begin
            superpage_entries_0_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_0_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1440) begin
            superpage_entries_0_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_0_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1440) begin
            superpage_entries_0_data_0 <= _T_1438;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_0_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      superpage_entries_0_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_0) begin
          superpage_entries_0_valid_0 <= 1'h0;
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_1439) begin
              superpage_entries_0_valid_0 <= _GEN_67;
            end
          end
        end
      end else begin
        superpage_entries_0_valid_0 <= _GEN_862;
      end
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          superpage_entries_0_valid_0 <= _GEN_67;
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_level <= 2'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1456) begin
            superpage_entries_1_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1456) begin
            superpage_entries_1_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1456) begin
            superpage_entries_1_data_0 <= _T_1438;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      superpage_entries_1_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_1) begin
          superpage_entries_1_valid_0 <= 1'h0;
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_1439) begin
              superpage_entries_1_valid_0 <= _GEN_71;
            end
          end
        end
      end else begin
        superpage_entries_1_valid_0 <= _GEN_866;
      end
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          superpage_entries_1_valid_0 <= _GEN_71;
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_level <= 2'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1472) begin
            superpage_entries_2_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1472) begin
            superpage_entries_2_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1472) begin
            superpage_entries_2_data_0 <= _T_1438;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      superpage_entries_2_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_2) begin
          superpage_entries_2_valid_0 <= 1'h0;
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_1439) begin
              superpage_entries_2_valid_0 <= _GEN_75;
            end
          end
        end
      end else begin
        superpage_entries_2_valid_0 <= _GEN_870;
      end
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          superpage_entries_2_valid_0 <= _GEN_75;
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_level <= 2'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1488) begin
            superpage_entries_3_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_tag <= 27'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1488) begin
            superpage_entries_3_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          if (_T_1488) begin
            superpage_entries_3_data_0 <= _T_1438;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      superpage_entries_3_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_3) begin
          superpage_entries_3_valid_0 <= 1'h0;
        end else if (_T_1385) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_1439) begin
              superpage_entries_3_valid_0 <= _GEN_79;
            end
          end
        end
      end else begin
        superpage_entries_3_valid_0 <= _GEN_874;
      end
    end else if (_T_1385) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_1439) begin
          superpage_entries_3_valid_0 <= _GEN_79;
        end
      end
    end
    if (metaReset) begin
      special_entry_level <= 2'h0;
    end else if (_T_1385) begin
      if (~io_ptw_resp_bits_homogeneous) begin
        special_entry_level <= io_ptw_resp_bits_level;
      end
    end
    if (metaReset) begin
      special_entry_tag <= 27'h0;
    end else if (_T_1385) begin
      if (~io_ptw_resp_bits_homogeneous) begin
        special_entry_tag <= r_refill_tag;
      end
    end
    if (metaReset) begin
      special_entry_data_0 <= 34'h0;
    end else if (_T_1385) begin
      if (~io_ptw_resp_bits_homogeneous) begin
        special_entry_data_0 <= _T_1438;
      end
    end
    if (metaReset) begin
      special_entry_valid_0 <= 1'h0;
    end else if (_T_4530) begin
      special_entry_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_994) begin
          special_entry_valid_0 <= 1'h0;
        end else if (_T_1385) begin
          special_entry_valid_0 <= _GEN_355;
        end
      end else begin
        special_entry_valid_0 <= _GEN_878;
      end
    end else if (_T_1385) begin
      special_entry_valid_0 <= _GEN_355;
    end
    if (metaReset) begin
      state <= 2'h0;
    end else if (reset) begin
      state <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      state <= 2'h0;
    end else if (_T_2941) begin
      state <= 2'h3;
    end else if (io_ptw_resp_valid) begin
      state <= 2'h0;
    end else if (_T_2941) begin
      state <= 2'h3;
    end else if (_T_324) begin
      if (io_kill) begin
        state <= 2'h0;
      end else if (io_ptw_req_ready) begin
        if (io_sfence_valid) begin
          state <= 2'h3;
        end else begin
          state <= 2'h2;
        end
      end else if (io_sfence_valid) begin
        state <= 2'h0;
      end else if (_T_2809) begin
        state <= 2'h1;
      end
    end else if (_T_2809) begin
      state <= 2'h1;
    end
    if (metaReset) begin
      r_refill_tag <= 27'h0;
    end else if (_T_2809) begin
      r_refill_tag <= vpn;
    end
    if (metaReset) begin
      r_superpage_repl_addr <= 2'h0;
    end else if (_T_2809) begin
      if (_T_2830) begin
        r_superpage_repl_addr <= _T_2824[1:0];
      end else if (_T_2832) begin
        r_superpage_repl_addr <= 2'h0;
      end else if (_T_2833) begin
        r_superpage_repl_addr <= 2'h1;
      end else if (_T_2834) begin
        r_superpage_repl_addr <= 2'h2;
      end else begin
        r_superpage_repl_addr <= 2'h3;
      end
    end
    if (metaReset) begin
      r_sectored_repl_addr <= 3'h0;
    end else if (_T_2809) begin
      if (_T_2895) begin
        r_sectored_repl_addr <= _T_2861[2:0];
      end else if (_T_2897) begin
        r_sectored_repl_addr <= 3'h0;
      end else if (_T_2898) begin
        r_sectored_repl_addr <= 3'h1;
      end else if (_T_2899) begin
        r_sectored_repl_addr <= 3'h2;
      end else if (_T_2900) begin
        r_sectored_repl_addr <= 3'h3;
      end else if (_T_2901) begin
        r_sectored_repl_addr <= 3'h4;
      end else if (_T_2902) begin
        r_sectored_repl_addr <= 3'h5;
      end else if (_T_2903) begin
        r_sectored_repl_addr <= 3'h6;
      end else begin
        r_sectored_repl_addr <= 3'h7;
      end
    end
    if (metaReset) begin
      r_sectored_hit_addr <= 3'h0;
    end else if (_T_2809) begin
      r_sectored_hit_addr <= _T_2582;
    end
    if (metaReset) begin
      r_sectored_hit <= 1'h0;
    end else if (_T_2809) begin
      r_sectored_hit <= _T_2564;
    end
    if (metaReset) begin
      vpoffset_cfg_value <= 27'h0;
    end else if (reset) begin
      vpoffset_cfg_value <= 27'h0;
    end else begin
      vpoffset_cfg_value <= io_ptw_vpoffset_bits_value;
    end
    if (metaReset) begin
      requestedVPN <= 27'h0;
    end else if (io_ptw_req_bits_valid) begin
      requestedVPN <= io_ptw_req_bits_bits_addr;
    end
    if (metaReset) begin
      _T_2554 <= 7'h0;
    end else if (_T_2557) begin
      if (_T_2564) begin
        _T_2554 <= _T_2609[7:1];
      end
    end
    if (metaReset) begin
      _T_2556 <= 3'h0;
    end else if (_T_2557) begin
      if (_T_2614) begin
        _T_2556 <= _T_2641[3:1];
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_sfence_valid & ~_T_2949) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TLB.scala:414 assert(!io.sfence.bits.rs1 || (io.sfence.bits.addr >> pgIdxBits) === vpn)\n"); // @[TLB.scala 414:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_sfence_valid & ~_T_2949) begin
          $fatal; // @[TLB.scala 414:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    TLB_1_state <= TLB_1_xor0;
    if (!(TLB_1_cov_read_data)) begin
      TLB_1_covSum <= TLB_1_covSum + 1'h1;
    end
    if (metaReset) begin
      TLB_1_metaAssert <= 1'h0;
    end else begin
      TLB_1_metaAssert <= TLB_1_metaAssert | TLB_1_or0;
    end
  end
  always @(posedge clock) begin
    if(TLB_1_cov_write_en & TLB_1_cov_write_mask) begin
      TLB_1_cov[TLB_1_cov_write_addr] <= TLB_1_cov_write_data; // @[Coverage map for TLB_1]
    end
  end
endmodule
module BTB(
  input         clock,
  input         reset,
  input  [38:0] io_req_bits_addr,
  output        io_resp_valid,
  output        io_resp_bits_taken,
  output        io_resp_bits_bridx,
  output [38:0] io_resp_bits_target,
  output [4:0]  io_resp_bits_entry,
  output [7:0]  io_resp_bits_bht_history,
  output        io_resp_bits_bht_value,
  input         io_btb_update_valid,
  input  [4:0]  io_btb_update_bits_prediction_entry,
  input  [38:0] io_btb_update_bits_pc,
  input         io_btb_update_bits_isValid,
  input  [38:0] io_btb_update_bits_br_pc,
  input  [1:0]  io_btb_update_bits_cfiType,
  input         io_bht_update_valid,
  input  [7:0]  io_bht_update_bits_prediction_history,
  input  [38:0] io_bht_update_bits_pc,
  input         io_bht_update_bits_branch,
  input         io_bht_update_bits_taken,
  input         io_bht_update_bits_mispredict,
  input         io_bht_advance_valid,
  input         io_bht_advance_bits_bht_value,
  input         io_ras_update_valid,
  input  [1:0]  io_ras_update_bits_cfiType,
  input  [38:0] io_ras_update_bits_returnAddr,
  output        io_ras_head_valid,
  output [38:0] io_ras_head_bits,
  input         io_flush,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg  _T_1161 [0:511]; // @[BTB.scala 113:26]
  reg [31:0] _RAND_0;
  wire  _T_1161__T_1232_data; // @[BTB.scala 113:26]
  wire [8:0] _T_1161__T_1232_addr; // @[BTB.scala 113:26]
  wire  _T_1161__T_1245_data; // @[BTB.scala 113:26]
  wire [8:0] _T_1161__T_1245_addr; // @[BTB.scala 113:26]
  wire  _T_1161__T_1245_mask; // @[BTB.scala 113:26]
  wire  _T_1161__T_1245_en; // @[BTB.scala 113:26]
  reg [12:0] idxs_0; // @[BTB.scala 188:17]
  reg [31:0] _RAND_1;
  reg [12:0] idxs_1; // @[BTB.scala 188:17]
  reg [31:0] _RAND_2;
  reg [12:0] idxs_2; // @[BTB.scala 188:17]
  reg [31:0] _RAND_3;
  reg [12:0] idxs_3; // @[BTB.scala 188:17]
  reg [31:0] _RAND_4;
  reg [12:0] idxs_4; // @[BTB.scala 188:17]
  reg [31:0] _RAND_5;
  reg [12:0] idxs_5; // @[BTB.scala 188:17]
  reg [31:0] _RAND_6;
  reg [12:0] idxs_6; // @[BTB.scala 188:17]
  reg [31:0] _RAND_7;
  reg [12:0] idxs_7; // @[BTB.scala 188:17]
  reg [31:0] _RAND_8;
  reg [12:0] idxs_8; // @[BTB.scala 188:17]
  reg [31:0] _RAND_9;
  reg [12:0] idxs_9; // @[BTB.scala 188:17]
  reg [31:0] _RAND_10;
  reg [12:0] idxs_10; // @[BTB.scala 188:17]
  reg [31:0] _RAND_11;
  reg [12:0] idxs_11; // @[BTB.scala 188:17]
  reg [31:0] _RAND_12;
  reg [12:0] idxs_12; // @[BTB.scala 188:17]
  reg [31:0] _RAND_13;
  reg [12:0] idxs_13; // @[BTB.scala 188:17]
  reg [31:0] _RAND_14;
  reg [12:0] idxs_14; // @[BTB.scala 188:17]
  reg [31:0] _RAND_15;
  reg [12:0] idxs_15; // @[BTB.scala 188:17]
  reg [31:0] _RAND_16;
  reg [12:0] idxs_16; // @[BTB.scala 188:17]
  reg [31:0] _RAND_17;
  reg [12:0] idxs_17; // @[BTB.scala 188:17]
  reg [31:0] _RAND_18;
  reg [12:0] idxs_18; // @[BTB.scala 188:17]
  reg [31:0] _RAND_19;
  reg [12:0] idxs_19; // @[BTB.scala 188:17]
  reg [31:0] _RAND_20;
  reg [12:0] idxs_20; // @[BTB.scala 188:17]
  reg [31:0] _RAND_21;
  reg [12:0] idxs_21; // @[BTB.scala 188:17]
  reg [31:0] _RAND_22;
  reg [12:0] idxs_22; // @[BTB.scala 188:17]
  reg [31:0] _RAND_23;
  reg [12:0] idxs_23; // @[BTB.scala 188:17]
  reg [31:0] _RAND_24;
  reg [12:0] idxs_24; // @[BTB.scala 188:17]
  reg [31:0] _RAND_25;
  reg [12:0] idxs_25; // @[BTB.scala 188:17]
  reg [31:0] _RAND_26;
  reg [12:0] idxs_26; // @[BTB.scala 188:17]
  reg [31:0] _RAND_27;
  reg [12:0] idxs_27; // @[BTB.scala 188:17]
  reg [31:0] _RAND_28;
  reg [2:0] idxPages_0; // @[BTB.scala 189:21]
  reg [31:0] _RAND_29;
  reg [2:0] idxPages_1; // @[BTB.scala 189:21]
  reg [31:0] _RAND_30;
  reg [2:0] idxPages_2; // @[BTB.scala 189:21]
  reg [31:0] _RAND_31;
  reg [2:0] idxPages_3; // @[BTB.scala 189:21]
  reg [31:0] _RAND_32;
  reg [2:0] idxPages_4; // @[BTB.scala 189:21]
  reg [31:0] _RAND_33;
  reg [2:0] idxPages_5; // @[BTB.scala 189:21]
  reg [31:0] _RAND_34;
  reg [2:0] idxPages_6; // @[BTB.scala 189:21]
  reg [31:0] _RAND_35;
  reg [2:0] idxPages_7; // @[BTB.scala 189:21]
  reg [31:0] _RAND_36;
  reg [2:0] idxPages_8; // @[BTB.scala 189:21]
  reg [31:0] _RAND_37;
  reg [2:0] idxPages_9; // @[BTB.scala 189:21]
  reg [31:0] _RAND_38;
  reg [2:0] idxPages_10; // @[BTB.scala 189:21]
  reg [31:0] _RAND_39;
  reg [2:0] idxPages_11; // @[BTB.scala 189:21]
  reg [31:0] _RAND_40;
  reg [2:0] idxPages_12; // @[BTB.scala 189:21]
  reg [31:0] _RAND_41;
  reg [2:0] idxPages_13; // @[BTB.scala 189:21]
  reg [31:0] _RAND_42;
  reg [2:0] idxPages_14; // @[BTB.scala 189:21]
  reg [31:0] _RAND_43;
  reg [2:0] idxPages_15; // @[BTB.scala 189:21]
  reg [31:0] _RAND_44;
  reg [2:0] idxPages_16; // @[BTB.scala 189:21]
  reg [31:0] _RAND_45;
  reg [2:0] idxPages_17; // @[BTB.scala 189:21]
  reg [31:0] _RAND_46;
  reg [2:0] idxPages_18; // @[BTB.scala 189:21]
  reg [31:0] _RAND_47;
  reg [2:0] idxPages_19; // @[BTB.scala 189:21]
  reg [31:0] _RAND_48;
  reg [2:0] idxPages_20; // @[BTB.scala 189:21]
  reg [31:0] _RAND_49;
  reg [2:0] idxPages_21; // @[BTB.scala 189:21]
  reg [31:0] _RAND_50;
  reg [2:0] idxPages_22; // @[BTB.scala 189:21]
  reg [31:0] _RAND_51;
  reg [2:0] idxPages_23; // @[BTB.scala 189:21]
  reg [31:0] _RAND_52;
  reg [2:0] idxPages_24; // @[BTB.scala 189:21]
  reg [31:0] _RAND_53;
  reg [2:0] idxPages_25; // @[BTB.scala 189:21]
  reg [31:0] _RAND_54;
  reg [2:0] idxPages_26; // @[BTB.scala 189:21]
  reg [31:0] _RAND_55;
  reg [2:0] idxPages_27; // @[BTB.scala 189:21]
  reg [31:0] _RAND_56;
  reg [12:0] tgts_0; // @[BTB.scala 190:17]
  reg [31:0] _RAND_57;
  reg [12:0] tgts_1; // @[BTB.scala 190:17]
  reg [31:0] _RAND_58;
  reg [12:0] tgts_2; // @[BTB.scala 190:17]
  reg [31:0] _RAND_59;
  reg [12:0] tgts_3; // @[BTB.scala 190:17]
  reg [31:0] _RAND_60;
  reg [12:0] tgts_4; // @[BTB.scala 190:17]
  reg [31:0] _RAND_61;
  reg [12:0] tgts_5; // @[BTB.scala 190:17]
  reg [31:0] _RAND_62;
  reg [12:0] tgts_6; // @[BTB.scala 190:17]
  reg [31:0] _RAND_63;
  reg [12:0] tgts_7; // @[BTB.scala 190:17]
  reg [31:0] _RAND_64;
  reg [12:0] tgts_8; // @[BTB.scala 190:17]
  reg [31:0] _RAND_65;
  reg [12:0] tgts_9; // @[BTB.scala 190:17]
  reg [31:0] _RAND_66;
  reg [12:0] tgts_10; // @[BTB.scala 190:17]
  reg [31:0] _RAND_67;
  reg [12:0] tgts_11; // @[BTB.scala 190:17]
  reg [31:0] _RAND_68;
  reg [12:0] tgts_12; // @[BTB.scala 190:17]
  reg [31:0] _RAND_69;
  reg [12:0] tgts_13; // @[BTB.scala 190:17]
  reg [31:0] _RAND_70;
  reg [12:0] tgts_14; // @[BTB.scala 190:17]
  reg [31:0] _RAND_71;
  reg [12:0] tgts_15; // @[BTB.scala 190:17]
  reg [31:0] _RAND_72;
  reg [12:0] tgts_16; // @[BTB.scala 190:17]
  reg [31:0] _RAND_73;
  reg [12:0] tgts_17; // @[BTB.scala 190:17]
  reg [31:0] _RAND_74;
  reg [12:0] tgts_18; // @[BTB.scala 190:17]
  reg [31:0] _RAND_75;
  reg [12:0] tgts_19; // @[BTB.scala 190:17]
  reg [31:0] _RAND_76;
  reg [12:0] tgts_20; // @[BTB.scala 190:17]
  reg [31:0] _RAND_77;
  reg [12:0] tgts_21; // @[BTB.scala 190:17]
  reg [31:0] _RAND_78;
  reg [12:0] tgts_22; // @[BTB.scala 190:17]
  reg [31:0] _RAND_79;
  reg [12:0] tgts_23; // @[BTB.scala 190:17]
  reg [31:0] _RAND_80;
  reg [12:0] tgts_24; // @[BTB.scala 190:17]
  reg [31:0] _RAND_81;
  reg [12:0] tgts_25; // @[BTB.scala 190:17]
  reg [31:0] _RAND_82;
  reg [12:0] tgts_26; // @[BTB.scala 190:17]
  reg [31:0] _RAND_83;
  reg [12:0] tgts_27; // @[BTB.scala 190:17]
  reg [31:0] _RAND_84;
  reg [2:0] tgtPages_0; // @[BTB.scala 191:21]
  reg [31:0] _RAND_85;
  reg [2:0] tgtPages_1; // @[BTB.scala 191:21]
  reg [31:0] _RAND_86;
  reg [2:0] tgtPages_2; // @[BTB.scala 191:21]
  reg [31:0] _RAND_87;
  reg [2:0] tgtPages_3; // @[BTB.scala 191:21]
  reg [31:0] _RAND_88;
  reg [2:0] tgtPages_4; // @[BTB.scala 191:21]
  reg [31:0] _RAND_89;
  reg [2:0] tgtPages_5; // @[BTB.scala 191:21]
  reg [31:0] _RAND_90;
  reg [2:0] tgtPages_6; // @[BTB.scala 191:21]
  reg [31:0] _RAND_91;
  reg [2:0] tgtPages_7; // @[BTB.scala 191:21]
  reg [31:0] _RAND_92;
  reg [2:0] tgtPages_8; // @[BTB.scala 191:21]
  reg [31:0] _RAND_93;
  reg [2:0] tgtPages_9; // @[BTB.scala 191:21]
  reg [31:0] _RAND_94;
  reg [2:0] tgtPages_10; // @[BTB.scala 191:21]
  reg [31:0] _RAND_95;
  reg [2:0] tgtPages_11; // @[BTB.scala 191:21]
  reg [31:0] _RAND_96;
  reg [2:0] tgtPages_12; // @[BTB.scala 191:21]
  reg [31:0] _RAND_97;
  reg [2:0] tgtPages_13; // @[BTB.scala 191:21]
  reg [31:0] _RAND_98;
  reg [2:0] tgtPages_14; // @[BTB.scala 191:21]
  reg [31:0] _RAND_99;
  reg [2:0] tgtPages_15; // @[BTB.scala 191:21]
  reg [31:0] _RAND_100;
  reg [2:0] tgtPages_16; // @[BTB.scala 191:21]
  reg [31:0] _RAND_101;
  reg [2:0] tgtPages_17; // @[BTB.scala 191:21]
  reg [31:0] _RAND_102;
  reg [2:0] tgtPages_18; // @[BTB.scala 191:21]
  reg [31:0] _RAND_103;
  reg [2:0] tgtPages_19; // @[BTB.scala 191:21]
  reg [31:0] _RAND_104;
  reg [2:0] tgtPages_20; // @[BTB.scala 191:21]
  reg [31:0] _RAND_105;
  reg [2:0] tgtPages_21; // @[BTB.scala 191:21]
  reg [31:0] _RAND_106;
  reg [2:0] tgtPages_22; // @[BTB.scala 191:21]
  reg [31:0] _RAND_107;
  reg [2:0] tgtPages_23; // @[BTB.scala 191:21]
  reg [31:0] _RAND_108;
  reg [2:0] tgtPages_24; // @[BTB.scala 191:21]
  reg [31:0] _RAND_109;
  reg [2:0] tgtPages_25; // @[BTB.scala 191:21]
  reg [31:0] _RAND_110;
  reg [2:0] tgtPages_26; // @[BTB.scala 191:21]
  reg [31:0] _RAND_111;
  reg [2:0] tgtPages_27; // @[BTB.scala 191:21]
  reg [31:0] _RAND_112;
  reg [24:0] pages_0; // @[BTB.scala 192:18]
  reg [31:0] _RAND_113;
  reg [24:0] pages_1; // @[BTB.scala 192:18]
  reg [31:0] _RAND_114;
  reg [24:0] pages_2; // @[BTB.scala 192:18]
  reg [31:0] _RAND_115;
  reg [24:0] pages_3; // @[BTB.scala 192:18]
  reg [31:0] _RAND_116;
  reg [24:0] pages_4; // @[BTB.scala 192:18]
  reg [31:0] _RAND_117;
  reg [24:0] pages_5; // @[BTB.scala 192:18]
  reg [31:0] _RAND_118;
  reg [5:0] pageValid; // @[BTB.scala 193:22]
  reg [31:0] _RAND_119;
  reg [27:0] isValid; // @[BTB.scala 195:20]
  reg [31:0] _RAND_120;
  reg [1:0] cfiType_0; // @[BTB.scala 196:20]
  reg [31:0] _RAND_121;
  reg [1:0] cfiType_1; // @[BTB.scala 196:20]
  reg [31:0] _RAND_122;
  reg [1:0] cfiType_2; // @[BTB.scala 196:20]
  reg [31:0] _RAND_123;
  reg [1:0] cfiType_3; // @[BTB.scala 196:20]
  reg [31:0] _RAND_124;
  reg [1:0] cfiType_4; // @[BTB.scala 196:20]
  reg [31:0] _RAND_125;
  reg [1:0] cfiType_5; // @[BTB.scala 196:20]
  reg [31:0] _RAND_126;
  reg [1:0] cfiType_6; // @[BTB.scala 196:20]
  reg [31:0] _RAND_127;
  reg [1:0] cfiType_7; // @[BTB.scala 196:20]
  reg [31:0] _RAND_128;
  reg [1:0] cfiType_8; // @[BTB.scala 196:20]
  reg [31:0] _RAND_129;
  reg [1:0] cfiType_9; // @[BTB.scala 196:20]
  reg [31:0] _RAND_130;
  reg [1:0] cfiType_10; // @[BTB.scala 196:20]
  reg [31:0] _RAND_131;
  reg [1:0] cfiType_11; // @[BTB.scala 196:20]
  reg [31:0] _RAND_132;
  reg [1:0] cfiType_12; // @[BTB.scala 196:20]
  reg [31:0] _RAND_133;
  reg [1:0] cfiType_13; // @[BTB.scala 196:20]
  reg [31:0] _RAND_134;
  reg [1:0] cfiType_14; // @[BTB.scala 196:20]
  reg [31:0] _RAND_135;
  reg [1:0] cfiType_15; // @[BTB.scala 196:20]
  reg [31:0] _RAND_136;
  reg [1:0] cfiType_16; // @[BTB.scala 196:20]
  reg [31:0] _RAND_137;
  reg [1:0] cfiType_17; // @[BTB.scala 196:20]
  reg [31:0] _RAND_138;
  reg [1:0] cfiType_18; // @[BTB.scala 196:20]
  reg [31:0] _RAND_139;
  reg [1:0] cfiType_19; // @[BTB.scala 196:20]
  reg [31:0] _RAND_140;
  reg [1:0] cfiType_20; // @[BTB.scala 196:20]
  reg [31:0] _RAND_141;
  reg [1:0] cfiType_21; // @[BTB.scala 196:20]
  reg [31:0] _RAND_142;
  reg [1:0] cfiType_22; // @[BTB.scala 196:20]
  reg [31:0] _RAND_143;
  reg [1:0] cfiType_23; // @[BTB.scala 196:20]
  reg [31:0] _RAND_144;
  reg [1:0] cfiType_24; // @[BTB.scala 196:20]
  reg [31:0] _RAND_145;
  reg [1:0] cfiType_25; // @[BTB.scala 196:20]
  reg [31:0] _RAND_146;
  reg [1:0] cfiType_26; // @[BTB.scala 196:20]
  reg [31:0] _RAND_147;
  reg [1:0] cfiType_27; // @[BTB.scala 196:20]
  reg [31:0] _RAND_148;
  reg  brIdx_0; // @[BTB.scala 197:18]
  reg [31:0] _RAND_149;
  reg  brIdx_1; // @[BTB.scala 197:18]
  reg [31:0] _RAND_150;
  reg  brIdx_2; // @[BTB.scala 197:18]
  reg [31:0] _RAND_151;
  reg  brIdx_3; // @[BTB.scala 197:18]
  reg [31:0] _RAND_152;
  reg  brIdx_4; // @[BTB.scala 197:18]
  reg [31:0] _RAND_153;
  reg  brIdx_5; // @[BTB.scala 197:18]
  reg [31:0] _RAND_154;
  reg  brIdx_6; // @[BTB.scala 197:18]
  reg [31:0] _RAND_155;
  reg  brIdx_7; // @[BTB.scala 197:18]
  reg [31:0] _RAND_156;
  reg  brIdx_8; // @[BTB.scala 197:18]
  reg [31:0] _RAND_157;
  reg  brIdx_9; // @[BTB.scala 197:18]
  reg [31:0] _RAND_158;
  reg  brIdx_10; // @[BTB.scala 197:18]
  reg [31:0] _RAND_159;
  reg  brIdx_11; // @[BTB.scala 197:18]
  reg [31:0] _RAND_160;
  reg  brIdx_12; // @[BTB.scala 197:18]
  reg [31:0] _RAND_161;
  reg  brIdx_13; // @[BTB.scala 197:18]
  reg [31:0] _RAND_162;
  reg  brIdx_14; // @[BTB.scala 197:18]
  reg [31:0] _RAND_163;
  reg  brIdx_15; // @[BTB.scala 197:18]
  reg [31:0] _RAND_164;
  reg  brIdx_16; // @[BTB.scala 197:18]
  reg [31:0] _RAND_165;
  reg  brIdx_17; // @[BTB.scala 197:18]
  reg [31:0] _RAND_166;
  reg  brIdx_18; // @[BTB.scala 197:18]
  reg [31:0] _RAND_167;
  reg  brIdx_19; // @[BTB.scala 197:18]
  reg [31:0] _RAND_168;
  reg  brIdx_20; // @[BTB.scala 197:18]
  reg [31:0] _RAND_169;
  reg  brIdx_21; // @[BTB.scala 197:18]
  reg [31:0] _RAND_170;
  reg  brIdx_22; // @[BTB.scala 197:18]
  reg [31:0] _RAND_171;
  reg  brIdx_23; // @[BTB.scala 197:18]
  reg [31:0] _RAND_172;
  reg  brIdx_24; // @[BTB.scala 197:18]
  reg [31:0] _RAND_173;
  reg  brIdx_25; // @[BTB.scala 197:18]
  reg [31:0] _RAND_174;
  reg  brIdx_26; // @[BTB.scala 197:18]
  reg [31:0] _RAND_175;
  reg  brIdx_27; // @[BTB.scala 197:18]
  reg [31:0] _RAND_176;
  reg  r_btb_update_valid; // @[Valid.scala 48:22]
  reg [31:0] _RAND_177;
  reg [4:0] r_btb_update_bits_prediction_entry; // @[Reg.scala 11:16]
  reg [31:0] _RAND_178;
  reg [38:0] r_btb_update_bits_pc; // @[Reg.scala 11:16]
  reg [63:0] _RAND_179;
  reg  r_btb_update_bits_isValid; // @[Reg.scala 11:16]
  reg [31:0] _RAND_180;
  reg [38:0] r_btb_update_bits_br_pc; // @[Reg.scala 11:16]
  reg [63:0] _RAND_181;
  reg [1:0] r_btb_update_bits_cfiType; // @[Reg.scala 11:16]
  reg [31:0] _RAND_182;
  wire  _T_249; // @[BTB.scala 202:29]
  wire  _T_250; // @[BTB.scala 202:29]
  wire  _T_251; // @[BTB.scala 202:29]
  wire  _T_252; // @[BTB.scala 202:29]
  wire  _T_253; // @[BTB.scala 202:29]
  wire  _T_254; // @[BTB.scala 202:29]
  wire [5:0] _T_259; // @[Cat.scala 30:58]
  wire [5:0] pageHit; // @[BTB.scala 202:15]
  wire  _T_261; // @[BTB.scala 206:16]
  wire  _T_262; // @[BTB.scala 206:16]
  wire  _T_263; // @[BTB.scala 206:16]
  wire  _T_264; // @[BTB.scala 206:16]
  wire  _T_265; // @[BTB.scala 206:16]
  wire  _T_266; // @[BTB.scala 206:16]
  wire  _T_267; // @[BTB.scala 206:16]
  wire  _T_268; // @[BTB.scala 206:16]
  wire  _T_269; // @[BTB.scala 206:16]
  wire  _T_270; // @[BTB.scala 206:16]
  wire  _T_271; // @[BTB.scala 206:16]
  wire  _T_272; // @[BTB.scala 206:16]
  wire  _T_273; // @[BTB.scala 206:16]
  wire  _T_274; // @[BTB.scala 206:16]
  wire  _T_275; // @[BTB.scala 206:16]
  wire  _T_276; // @[BTB.scala 206:16]
  wire  _T_277; // @[BTB.scala 206:16]
  wire  _T_278; // @[BTB.scala 206:16]
  wire  _T_279; // @[BTB.scala 206:16]
  wire  _T_280; // @[BTB.scala 206:16]
  wire  _T_281; // @[BTB.scala 206:16]
  wire  _T_282; // @[BTB.scala 206:16]
  wire  _T_283; // @[BTB.scala 206:16]
  wire  _T_284; // @[BTB.scala 206:16]
  wire  _T_285; // @[BTB.scala 206:16]
  wire  _T_286; // @[BTB.scala 206:16]
  wire  _T_287; // @[BTB.scala 206:16]
  wire  _T_288; // @[BTB.scala 206:16]
  wire [6:0] _T_294; // @[Cat.scala 30:58]
  wire [13:0] _T_301; // @[Cat.scala 30:58]
  wire [6:0] _T_307; // @[Cat.scala 30:58]
  wire [27:0] _T_315; // @[Cat.scala 30:58]
  wire [27:0] idxHit; // @[BTB.scala 206:32]
  wire  _T_317; // @[BTB.scala 202:29]
  wire  _T_318; // @[BTB.scala 202:29]
  wire  _T_319; // @[BTB.scala 202:29]
  wire  _T_320; // @[BTB.scala 202:29]
  wire  _T_321; // @[BTB.scala 202:29]
  wire  _T_322; // @[BTB.scala 202:29]
  wire [5:0] _T_327; // @[Cat.scala 30:58]
  wire [5:0] updatePageHit; // @[BTB.scala 202:15]
  wire  updateHit; // @[BTB.scala 220:48]
  wire  useUpdatePageHit; // @[BTB.scala 222:40]
  wire  usePageHit; // @[BTB.scala 223:28]
  wire  doIdxPageRepl; // @[BTB.scala 224:23]
  reg [2:0] nextPageRepl; // @[BTB.scala 225:25]
  reg [31:0] _RAND_183;
  wire [5:0] _T_331; // @[Cat.scala 30:58]
  wire [7:0] _T_332; // @[OneHot.scala 45:35]
  wire [7:0] _T_333; // @[BTB.scala 226:70]
  wire [7:0] _GEN_432; // @[BTB.scala 226:65]
  wire [7:0] idxPageRepl; // @[BTB.scala 226:65]
  wire [7:0] idxPageUpdateOH; // @[BTB.scala 227:28]
  wire  _T_336; // @[OneHot.scala 28:14]
  wire [3:0] _T_337; // @[OneHot.scala 28:28]
  wire  _T_340; // @[OneHot.scala 28:14]
  wire [1:0] _T_341; // @[OneHot.scala 28:28]
  wire [2:0] idxPageUpdate; // @[Cat.scala 30:58]
  wire [7:0] idxPageReplEn; // @[BTB.scala 229:26]
  wire  samePage; // @[BTB.scala 231:45]
  wire  doTgtPageRepl; // @[BTB.scala 232:33]
  wire [5:0] _T_350; // @[Cat.scala 30:58]
  wire [7:0] tgtPageRepl; // @[BTB.scala 233:24]
  wire [7:0] _T_351; // @[BTB.scala 234:45]
  wire [7:0] _GEN_433; // @[BTB.scala 234:40]
  wire [7:0] _T_352; // @[BTB.scala 234:40]
  wire  _T_355; // @[OneHot.scala 28:14]
  wire [3:0] _T_356; // @[OneHot.scala 28:28]
  wire  _T_359; // @[OneHot.scala 28:14]
  wire [1:0] _T_360; // @[OneHot.scala 28:28]
  wire [2:0] tgtPageUpdate; // @[Cat.scala 30:58]
  wire [7:0] tgtPageReplEn; // @[BTB.scala 235:26]
  wire  _T_363; // @[BTB.scala 237:46]
  wire  _T_364; // @[BTB.scala 237:28]
  wire  _T_365; // @[BTB.scala 238:30]
  wire [1:0] _T_366; // @[BTB.scala 239:40]
  wire [2:0] _GEN_434; // @[BTB.scala 239:29]
  wire [2:0] _T_368; // @[BTB.scala 239:29]
  wire  _T_369; // @[BTB.scala 240:30]
  reg [26:0] _T_373; // @[Replacement.scala 41:30]
  reg [31:0] _RAND_184;
  wire [27:0] _T_374; // @[Replacement.scala 57:31]
  wire [27:0] _T_378; // @[Replacement.scala 61:48]
  wire [1:0] _T_381; // @[Cat.scala 30:58]
  wire [5:0] _T_382; // @[Cat.scala 30:58]
  wire  _T_384; // @[Replacement.scala 60:70]
  wire [27:0] _T_385; // @[Replacement.scala 61:48]
  wire  _T_387; // @[Replacement.scala 61:32]
  wire [2:0] _T_388; // @[Cat.scala 30:58]
  wire [5:0] _T_389; // @[Cat.scala 30:58]
  wire  _T_391; // @[Replacement.scala 60:70]
  wire [27:0] _T_392; // @[Replacement.scala 61:48]
  wire  _T_394; // @[Replacement.scala 61:32]
  wire [3:0] _T_395; // @[Cat.scala 30:58]
  wire [5:0] _T_396; // @[Cat.scala 30:58]
  wire  _T_398; // @[Replacement.scala 60:70]
  wire [27:0] _T_399; // @[Replacement.scala 61:48]
  wire  _T_401; // @[Replacement.scala 61:32]
  wire [4:0] _T_402; // @[Cat.scala 30:58]
  wire [5:0] _T_403; // @[Cat.scala 30:58]
  wire  _T_405; // @[Replacement.scala 60:70]
  wire [27:0] _T_406; // @[Replacement.scala 61:48]
  wire  _T_408; // @[Replacement.scala 61:32]
  wire [5:0] _T_409; // @[Cat.scala 30:58]
  wire [4:0] waddr; // @[BTB.scala 244:18]
  reg  r_resp_valid; // @[Valid.scala 48:22]
  reg [31:0] _RAND_185;
  reg  r_resp_bits_taken; // @[Reg.scala 11:16]
  reg [31:0] _RAND_186;
  reg [4:0] r_resp_bits_entry; // @[Reg.scala 11:16]
  reg [31:0] _RAND_187;
  wire  _T_419; // @[BTB.scala 246:22]
  wire  _T_420; // @[BTB.scala 246:43]
  wire [4:0] _T_421; // @[BTB.scala 247:20]
  wire [27:0] _T_426; // @[Replacement.scala 50:37]
  wire [27:0] _T_428; // @[Replacement.scala 50:37]
  wire [27:0] _T_430; // @[Replacement.scala 50:37]
  wire [1:0] _T_431; // @[Cat.scala 30:58]
  wire [3:0] _T_434; // @[Replacement.scala 50:37]
  wire [27:0] _GEN_436; // @[Replacement.scala 50:37]
  wire [27:0] _T_435; // @[Replacement.scala 50:37]
  wire [27:0] _T_437; // @[Replacement.scala 50:37]
  wire [27:0] _T_439; // @[Replacement.scala 50:37]
  wire [2:0] _T_440; // @[Cat.scala 30:58]
  wire [7:0] _T_443; // @[Replacement.scala 50:37]
  wire [27:0] _GEN_438; // @[Replacement.scala 50:37]
  wire [27:0] _T_444; // @[Replacement.scala 50:37]
  wire [27:0] _T_446; // @[Replacement.scala 50:37]
  wire [27:0] _T_448; // @[Replacement.scala 50:37]
  wire [3:0] _T_449; // @[Cat.scala 30:58]
  wire [15:0] _T_452; // @[Replacement.scala 50:37]
  wire [27:0] _GEN_440; // @[Replacement.scala 50:37]
  wire [27:0] _T_453; // @[Replacement.scala 50:37]
  wire [27:0] _T_455; // @[Replacement.scala 50:37]
  wire [27:0] _T_457; // @[Replacement.scala 50:37]
  wire [4:0] _T_458; // @[Cat.scala 30:58]
  wire [31:0] _T_461; // @[Replacement.scala 50:37]
  wire [31:0] _GEN_442; // @[Replacement.scala 50:37]
  wire [31:0] _T_462; // @[Replacement.scala 50:37]
  wire [31:0] _GEN_443; // @[Replacement.scala 50:37]
  wire [31:0] _T_464; // @[Replacement.scala 50:37]
  wire [31:0] _T_466; // @[Replacement.scala 50:37]
  wire [31:0] _T_469; // @[OneHot.scala 45:35]
  wire [3:0] _T_475; // @[BTB.scala 254:38]
  wire [31:0] _GEN_444; // @[BTB.scala 257:55]
  wire [31:0] _T_478; // @[BTB.scala 257:55]
  wire [31:0] _T_480; // @[BTB.scala 257:71]
  wire [31:0] _T_481; // @[BTB.scala 257:19]
  wire [7:0] _T_486; // @[BTB.scala 268:24]
  wire [7:0] _T_493; // @[BTB.scala 270:24]
  wire [7:0] _GEN_446; // @[BTB.scala 272:28]
  wire [7:0] _T_500; // @[BTB.scala 272:28]
  wire [7:0] _T_501; // @[BTB.scala 272:44]
  wire [31:0] _GEN_338; // @[BTB.scala 250:29]
  wire [7:0] _GEN_373; // @[BTB.scala 250:29]
  wire [6:0] _T_502; // @[BTB.scala 275:29]
  wire [2:0] _T_532; // @[Mux.scala 19:72]
  wire [2:0] _T_533; // @[Mux.scala 19:72]
  wire [2:0] _T_534; // @[Mux.scala 19:72]
  wire [2:0] _T_535; // @[Mux.scala 19:72]
  wire [2:0] _T_536; // @[Mux.scala 19:72]
  wire [2:0] _T_537; // @[Mux.scala 19:72]
  wire [2:0] _T_538; // @[Mux.scala 19:72]
  wire [2:0] _T_539; // @[Mux.scala 19:72]
  wire [2:0] _T_540; // @[Mux.scala 19:72]
  wire [2:0] _T_541; // @[Mux.scala 19:72]
  wire [2:0] _T_542; // @[Mux.scala 19:72]
  wire [2:0] _T_543; // @[Mux.scala 19:72]
  wire [2:0] _T_544; // @[Mux.scala 19:72]
  wire [2:0] _T_545; // @[Mux.scala 19:72]
  wire [2:0] _T_546; // @[Mux.scala 19:72]
  wire [2:0] _T_547; // @[Mux.scala 19:72]
  wire [2:0] _T_548; // @[Mux.scala 19:72]
  wire [2:0] _T_549; // @[Mux.scala 19:72]
  wire [2:0] _T_550; // @[Mux.scala 19:72]
  wire [2:0] _T_551; // @[Mux.scala 19:72]
  wire [2:0] _T_552; // @[Mux.scala 19:72]
  wire [2:0] _T_553; // @[Mux.scala 19:72]
  wire [2:0] _T_554; // @[Mux.scala 19:72]
  wire [2:0] _T_555; // @[Mux.scala 19:72]
  wire [2:0] _T_556; // @[Mux.scala 19:72]
  wire [2:0] _T_557; // @[Mux.scala 19:72]
  wire [2:0] _T_558; // @[Mux.scala 19:72]
  wire [2:0] _T_559; // @[Mux.scala 19:72]
  wire [2:0] _T_560; // @[Mux.scala 19:72]
  wire [2:0] _T_561; // @[Mux.scala 19:72]
  wire [2:0] _T_562; // @[Mux.scala 19:72]
  wire [2:0] _T_563; // @[Mux.scala 19:72]
  wire [2:0] _T_564; // @[Mux.scala 19:72]
  wire [2:0] _T_565; // @[Mux.scala 19:72]
  wire [2:0] _T_566; // @[Mux.scala 19:72]
  wire [2:0] _T_567; // @[Mux.scala 19:72]
  wire [2:0] _T_568; // @[Mux.scala 19:72]
  wire [2:0] _T_569; // @[Mux.scala 19:72]
  wire [2:0] _T_570; // @[Mux.scala 19:72]
  wire [2:0] _T_571; // @[Mux.scala 19:72]
  wire [2:0] _T_572; // @[Mux.scala 19:72]
  wire [2:0] _T_573; // @[Mux.scala 19:72]
  wire [2:0] _T_574; // @[Mux.scala 19:72]
  wire [2:0] _T_575; // @[Mux.scala 19:72]
  wire [2:0] _T_576; // @[Mux.scala 19:72]
  wire [2:0] _T_577; // @[Mux.scala 19:72]
  wire [2:0] _T_578; // @[Mux.scala 19:72]
  wire [2:0] _T_579; // @[Mux.scala 19:72]
  wire [2:0] _T_580; // @[Mux.scala 19:72]
  wire [2:0] _T_581; // @[Mux.scala 19:72]
  wire [2:0] _T_582; // @[Mux.scala 19:72]
  wire [2:0] _T_583; // @[Mux.scala 19:72]
  wire [2:0] _T_584; // @[Mux.scala 19:72]
  wire [2:0] _T_585; // @[Mux.scala 19:72]
  wire [2:0] _T_586; // @[Mux.scala 19:72]
  wire [6:0] _T_589; // @[BTB.scala 275:34]
  wire [2:0] _T_620; // @[Mux.scala 19:72]
  wire [2:0] _T_621; // @[Mux.scala 19:72]
  wire [2:0] _T_622; // @[Mux.scala 19:72]
  wire [2:0] _T_623; // @[Mux.scala 19:72]
  wire [2:0] _T_624; // @[Mux.scala 19:72]
  wire [2:0] _T_625; // @[Mux.scala 19:72]
  wire [2:0] _T_626; // @[Mux.scala 19:72]
  wire [2:0] _T_627; // @[Mux.scala 19:72]
  wire [2:0] _T_628; // @[Mux.scala 19:72]
  wire [2:0] _T_629; // @[Mux.scala 19:72]
  wire [2:0] _T_630; // @[Mux.scala 19:72]
  wire [2:0] _T_631; // @[Mux.scala 19:72]
  wire [2:0] _T_632; // @[Mux.scala 19:72]
  wire [2:0] _T_633; // @[Mux.scala 19:72]
  wire [2:0] _T_634; // @[Mux.scala 19:72]
  wire [2:0] _T_635; // @[Mux.scala 19:72]
  wire [2:0] _T_636; // @[Mux.scala 19:72]
  wire [2:0] _T_637; // @[Mux.scala 19:72]
  wire [2:0] _T_638; // @[Mux.scala 19:72]
  wire [2:0] _T_639; // @[Mux.scala 19:72]
  wire [2:0] _T_640; // @[Mux.scala 19:72]
  wire [2:0] _T_641; // @[Mux.scala 19:72]
  wire [2:0] _T_642; // @[Mux.scala 19:72]
  wire [2:0] _T_643; // @[Mux.scala 19:72]
  wire [2:0] _T_644; // @[Mux.scala 19:72]
  wire [2:0] _T_645; // @[Mux.scala 19:72]
  wire [2:0] _T_646; // @[Mux.scala 19:72]
  wire [2:0] _T_647; // @[Mux.scala 19:72]
  wire [2:0] _T_648; // @[Mux.scala 19:72]
  wire [2:0] _T_649; // @[Mux.scala 19:72]
  wire [2:0] _T_650; // @[Mux.scala 19:72]
  wire [2:0] _T_651; // @[Mux.scala 19:72]
  wire [2:0] _T_652; // @[Mux.scala 19:72]
  wire [2:0] _T_653; // @[Mux.scala 19:72]
  wire [2:0] _T_654; // @[Mux.scala 19:72]
  wire [2:0] _T_655; // @[Mux.scala 19:72]
  wire [2:0] _T_656; // @[Mux.scala 19:72]
  wire [2:0] _T_657; // @[Mux.scala 19:72]
  wire [2:0] _T_658; // @[Mux.scala 19:72]
  wire [2:0] _T_659; // @[Mux.scala 19:72]
  wire [2:0] _T_660; // @[Mux.scala 19:72]
  wire [2:0] _T_661; // @[Mux.scala 19:72]
  wire [2:0] _T_662; // @[Mux.scala 19:72]
  wire [2:0] _T_663; // @[Mux.scala 19:72]
  wire [2:0] _T_664; // @[Mux.scala 19:72]
  wire [2:0] _T_665; // @[Mux.scala 19:72]
  wire [2:0] _T_666; // @[Mux.scala 19:72]
  wire [2:0] _T_667; // @[Mux.scala 19:72]
  wire [2:0] _T_668; // @[Mux.scala 19:72]
  wire [2:0] _T_669; // @[Mux.scala 19:72]
  wire [2:0] _T_670; // @[Mux.scala 19:72]
  wire [2:0] _T_671; // @[Mux.scala 19:72]
  wire [2:0] _T_672; // @[Mux.scala 19:72]
  wire [2:0] _T_673; // @[Mux.scala 19:72]
  wire [2:0] _T_674; // @[Mux.scala 19:72]
  wire [12:0] _T_707; // @[Mux.scala 19:72]
  wire [12:0] _T_708; // @[Mux.scala 19:72]
  wire [12:0] _T_709; // @[Mux.scala 19:72]
  wire [12:0] _T_710; // @[Mux.scala 19:72]
  wire [12:0] _T_711; // @[Mux.scala 19:72]
  wire [12:0] _T_712; // @[Mux.scala 19:72]
  wire [12:0] _T_713; // @[Mux.scala 19:72]
  wire [12:0] _T_714; // @[Mux.scala 19:72]
  wire [12:0] _T_715; // @[Mux.scala 19:72]
  wire [12:0] _T_716; // @[Mux.scala 19:72]
  wire [12:0] _T_717; // @[Mux.scala 19:72]
  wire [12:0] _T_718; // @[Mux.scala 19:72]
  wire [12:0] _T_719; // @[Mux.scala 19:72]
  wire [12:0] _T_720; // @[Mux.scala 19:72]
  wire [12:0] _T_721; // @[Mux.scala 19:72]
  wire [12:0] _T_722; // @[Mux.scala 19:72]
  wire [12:0] _T_723; // @[Mux.scala 19:72]
  wire [12:0] _T_724; // @[Mux.scala 19:72]
  wire [12:0] _T_725; // @[Mux.scala 19:72]
  wire [12:0] _T_726; // @[Mux.scala 19:72]
  wire [12:0] _T_727; // @[Mux.scala 19:72]
  wire [12:0] _T_728; // @[Mux.scala 19:72]
  wire [12:0] _T_729; // @[Mux.scala 19:72]
  wire [12:0] _T_730; // @[Mux.scala 19:72]
  wire [12:0] _T_731; // @[Mux.scala 19:72]
  wire [12:0] _T_732; // @[Mux.scala 19:72]
  wire [12:0] _T_733; // @[Mux.scala 19:72]
  wire [12:0] _T_734; // @[Mux.scala 19:72]
  wire [12:0] _T_735; // @[Mux.scala 19:72]
  wire [12:0] _T_736; // @[Mux.scala 19:72]
  wire [12:0] _T_737; // @[Mux.scala 19:72]
  wire [12:0] _T_738; // @[Mux.scala 19:72]
  wire [12:0] _T_739; // @[Mux.scala 19:72]
  wire [12:0] _T_740; // @[Mux.scala 19:72]
  wire [12:0] _T_741; // @[Mux.scala 19:72]
  wire [12:0] _T_742; // @[Mux.scala 19:72]
  wire [12:0] _T_743; // @[Mux.scala 19:72]
  wire [12:0] _T_744; // @[Mux.scala 19:72]
  wire [12:0] _T_745; // @[Mux.scala 19:72]
  wire [12:0] _T_746; // @[Mux.scala 19:72]
  wire [12:0] _T_747; // @[Mux.scala 19:72]
  wire [12:0] _T_748; // @[Mux.scala 19:72]
  wire [12:0] _T_749; // @[Mux.scala 19:72]
  wire [12:0] _T_750; // @[Mux.scala 19:72]
  wire [12:0] _T_751; // @[Mux.scala 19:72]
  wire [12:0] _T_752; // @[Mux.scala 19:72]
  wire [12:0] _T_753; // @[Mux.scala 19:72]
  wire [12:0] _T_754; // @[Mux.scala 19:72]
  wire [12:0] _T_755; // @[Mux.scala 19:72]
  wire [12:0] _T_756; // @[Mux.scala 19:72]
  wire [12:0] _T_757; // @[Mux.scala 19:72]
  wire [12:0] _T_758; // @[Mux.scala 19:72]
  wire [12:0] _T_759; // @[Mux.scala 19:72]
  wire [12:0] _T_760; // @[Mux.scala 19:72]
  wire [12:0] _T_761; // @[Mux.scala 19:72]
  wire [13:0] _T_764; // @[BTB.scala 277:82]
  wire [24:0] _GEN_375; // @[Cat.scala 30:58]
  wire [24:0] _GEN_376; // @[Cat.scala 30:58]
  wire [24:0] _GEN_377; // @[Cat.scala 30:58]
  wire [24:0] _GEN_378; // @[Cat.scala 30:58]
  wire [24:0] _GEN_379; // @[Cat.scala 30:58]
  wire [38:0] _T_765; // @[Cat.scala 30:58]
  wire  _T_768; // @[OneHot.scala 28:14]
  wire [15:0] _GEN_447; // @[OneHot.scala 28:28]
  wire [15:0] _T_769; // @[OneHot.scala 28:28]
  wire  _T_772; // @[OneHot.scala 28:14]
  wire [7:0] _T_773; // @[OneHot.scala 28:28]
  wire  _T_776; // @[OneHot.scala 28:14]
  wire [3:0] _T_777; // @[OneHot.scala 28:28]
  wire  _T_780; // @[OneHot.scala 28:14]
  wire [1:0] _T_781; // @[OneHot.scala 28:28]
  wire [3:0] _T_785; // @[Cat.scala 30:58]
  wire  _T_816; // @[Mux.scala 19:72]
  wire  _T_817; // @[Mux.scala 19:72]
  wire  _T_818; // @[Mux.scala 19:72]
  wire  _T_819; // @[Mux.scala 19:72]
  wire  _T_820; // @[Mux.scala 19:72]
  wire  _T_821; // @[Mux.scala 19:72]
  wire  _T_822; // @[Mux.scala 19:72]
  wire  _T_823; // @[Mux.scala 19:72]
  wire  _T_824; // @[Mux.scala 19:72]
  wire  _T_825; // @[Mux.scala 19:72]
  wire  _T_826; // @[Mux.scala 19:72]
  wire  _T_827; // @[Mux.scala 19:72]
  wire  _T_828; // @[Mux.scala 19:72]
  wire  _T_829; // @[Mux.scala 19:72]
  wire  _T_830; // @[Mux.scala 19:72]
  wire  _T_831; // @[Mux.scala 19:72]
  wire  _T_832; // @[Mux.scala 19:72]
  wire  _T_833; // @[Mux.scala 19:72]
  wire  _T_834; // @[Mux.scala 19:72]
  wire  _T_835; // @[Mux.scala 19:72]
  wire  _T_836; // @[Mux.scala 19:72]
  wire  _T_837; // @[Mux.scala 19:72]
  wire  _T_838; // @[Mux.scala 19:72]
  wire  _T_839; // @[Mux.scala 19:72]
  wire  _T_840; // @[Mux.scala 19:72]
  wire  _T_841; // @[Mux.scala 19:72]
  wire  _T_842; // @[Mux.scala 19:72]
  wire  _T_843; // @[Mux.scala 19:72]
  wire  _T_844; // @[Mux.scala 19:72]
  wire  _T_845; // @[Mux.scala 19:72]
  wire  _T_846; // @[Mux.scala 19:72]
  wire  _T_847; // @[Mux.scala 19:72]
  wire  _T_848; // @[Mux.scala 19:72]
  wire  _T_849; // @[Mux.scala 19:72]
  wire  _T_850; // @[Mux.scala 19:72]
  wire  _T_851; // @[Mux.scala 19:72]
  wire  _T_852; // @[Mux.scala 19:72]
  wire  _T_853; // @[Mux.scala 19:72]
  wire  _T_854; // @[Mux.scala 19:72]
  wire  _T_855; // @[Mux.scala 19:72]
  wire  _T_856; // @[Mux.scala 19:72]
  wire  _T_857; // @[Mux.scala 19:72]
  wire  _T_858; // @[Mux.scala 19:72]
  wire  _T_859; // @[Mux.scala 19:72]
  wire  _T_860; // @[Mux.scala 19:72]
  wire  _T_861; // @[Mux.scala 19:72]
  wire  _T_862; // @[Mux.scala 19:72]
  wire  _T_863; // @[Mux.scala 19:72]
  wire  _T_864; // @[Mux.scala 19:72]
  wire  _T_865; // @[Mux.scala 19:72]
  wire  _T_866; // @[Mux.scala 19:72]
  wire  _T_867; // @[Mux.scala 19:72]
  wire  _T_868; // @[Mux.scala 19:72]
  wire  _T_869; // @[Mux.scala 19:72]
  wire  _T_977; // @[Misc.scala 187:16]
  wire  _T_979; // @[Misc.scala 187:61]
  wire  _T_981; // @[Misc.scala 187:16]
  wire  _T_983; // @[Misc.scala 187:61]
  wire  _T_984; // @[Misc.scala 187:49]
  wire  _T_991; // @[Misc.scala 187:16]
  wire  _T_993; // @[Misc.scala 187:61]
  wire  _T_1000; // @[Misc.scala 187:16]
  wire  _T_1002; // @[Misc.scala 187:61]
  wire  _T_1004; // @[Misc.scala 187:16]
  wire  _T_1005; // @[Misc.scala 187:37]
  wire  _T_1006; // @[Misc.scala 187:61]
  wire  _T_1007; // @[Misc.scala 187:49]
  wire  _T_1008; // @[Misc.scala 187:16]
  wire  _T_1009; // @[Misc.scala 187:37]
  wire  _T_1010; // @[Misc.scala 187:61]
  wire  _T_1011; // @[Misc.scala 187:49]
  wire  _T_1021; // @[Misc.scala 187:16]
  wire  _T_1023; // @[Misc.scala 187:61]
  wire  _T_1025; // @[Misc.scala 187:16]
  wire  _T_1027; // @[Misc.scala 187:61]
  wire  _T_1028; // @[Misc.scala 187:49]
  wire  _T_1035; // @[Misc.scala 187:16]
  wire  _T_1037; // @[Misc.scala 187:61]
  wire  _T_1044; // @[Misc.scala 187:16]
  wire  _T_1046; // @[Misc.scala 187:61]
  wire  _T_1048; // @[Misc.scala 187:16]
  wire  _T_1049; // @[Misc.scala 187:37]
  wire  _T_1050; // @[Misc.scala 187:61]
  wire  _T_1051; // @[Misc.scala 187:49]
  wire  _T_1052; // @[Misc.scala 187:16]
  wire  _T_1053; // @[Misc.scala 187:37]
  wire  _T_1054; // @[Misc.scala 187:61]
  wire  _T_1055; // @[Misc.scala 187:49]
  wire  _T_1056; // @[Misc.scala 187:16]
  wire  _T_1057; // @[Misc.scala 187:37]
  wire  _T_1058; // @[Misc.scala 187:61]
  wire  _T_1059; // @[Misc.scala 187:49]
  wire  _T_1070; // @[Misc.scala 187:16]
  wire  _T_1072; // @[Misc.scala 187:61]
  wire  _T_1074; // @[Misc.scala 187:16]
  wire  _T_1076; // @[Misc.scala 187:61]
  wire  _T_1077; // @[Misc.scala 187:49]
  wire  _T_1084; // @[Misc.scala 187:16]
  wire  _T_1086; // @[Misc.scala 187:61]
  wire  _T_1093; // @[Misc.scala 187:16]
  wire  _T_1095; // @[Misc.scala 187:61]
  wire  _T_1097; // @[Misc.scala 187:16]
  wire  _T_1098; // @[Misc.scala 187:37]
  wire  _T_1099; // @[Misc.scala 187:61]
  wire  _T_1100; // @[Misc.scala 187:49]
  wire  _T_1101; // @[Misc.scala 187:16]
  wire  _T_1102; // @[Misc.scala 187:37]
  wire  _T_1103; // @[Misc.scala 187:61]
  wire  _T_1104; // @[Misc.scala 187:49]
  wire  _T_1114; // @[Misc.scala 187:16]
  wire  _T_1116; // @[Misc.scala 187:61]
  wire  _T_1118; // @[Misc.scala 187:16]
  wire  _T_1120; // @[Misc.scala 187:61]
  wire  _T_1121; // @[Misc.scala 187:49]
  wire  _T_1128; // @[Misc.scala 187:16]
  wire  _T_1130; // @[Misc.scala 187:61]
  wire  _T_1137; // @[Misc.scala 187:16]
  wire  _T_1139; // @[Misc.scala 187:61]
  wire  _T_1141; // @[Misc.scala 187:16]
  wire  _T_1142; // @[Misc.scala 187:37]
  wire  _T_1143; // @[Misc.scala 187:61]
  wire  _T_1144; // @[Misc.scala 187:49]
  wire  _T_1145; // @[Misc.scala 187:16]
  wire  _T_1146; // @[Misc.scala 187:37]
  wire  _T_1147; // @[Misc.scala 187:61]
  wire  _T_1148; // @[Misc.scala 187:49]
  wire  _T_1149; // @[Misc.scala 187:16]
  wire  _T_1150; // @[Misc.scala 187:37]
  wire  _T_1151; // @[Misc.scala 187:61]
  wire  _T_1152; // @[Misc.scala 187:49]
  wire  _T_1154; // @[Misc.scala 187:37]
  wire  _T_1155; // @[Misc.scala 187:61]
  wire  _T_1156; // @[Misc.scala 187:49]
  wire [27:0] _T_1158; // @[BTB.scala 285:24]
  wire [31:0] _GEN_380; // @[BTB.scala 284:37]
  wire [31:0] _GEN_381; // @[BTB.scala 287:19]
  reg [7:0] _T_1163; // @[BTB.scala 114:20]
  reg [31:0] _RAND_188;
  wire  _T_1164; // @[BTB.scala 293:44]
  wire  _T_1165; // @[BTB.scala 293:44]
  wire  _T_1166; // @[BTB.scala 293:44]
  wire  _T_1167; // @[BTB.scala 293:44]
  wire  _T_1168; // @[BTB.scala 293:44]
  wire  _T_1169; // @[BTB.scala 293:44]
  wire  _T_1170; // @[BTB.scala 293:44]
  wire  _T_1171; // @[BTB.scala 293:44]
  wire  _T_1172; // @[BTB.scala 293:44]
  wire  _T_1173; // @[BTB.scala 293:44]
  wire  _T_1174; // @[BTB.scala 293:44]
  wire  _T_1175; // @[BTB.scala 293:44]
  wire  _T_1176; // @[BTB.scala 293:44]
  wire  _T_1177; // @[BTB.scala 293:44]
  wire  _T_1178; // @[BTB.scala 293:44]
  wire  _T_1179; // @[BTB.scala 293:44]
  wire  _T_1180; // @[BTB.scala 293:44]
  wire  _T_1181; // @[BTB.scala 293:44]
  wire  _T_1182; // @[BTB.scala 293:44]
  wire  _T_1183; // @[BTB.scala 293:44]
  wire  _T_1184; // @[BTB.scala 293:44]
  wire  _T_1185; // @[BTB.scala 293:44]
  wire  _T_1186; // @[BTB.scala 293:44]
  wire  _T_1187; // @[BTB.scala 293:44]
  wire  _T_1188; // @[BTB.scala 293:44]
  wire  _T_1189; // @[BTB.scala 293:44]
  wire  _T_1190; // @[BTB.scala 293:44]
  wire  _T_1191; // @[BTB.scala 293:44]
  wire [6:0] _T_1197; // @[Cat.scala 30:58]
  wire [13:0] _T_1204; // @[Cat.scala 30:58]
  wire [6:0] _T_1210; // @[Cat.scala 30:58]
  wire [27:0] _T_1218; // @[Cat.scala 30:58]
  wire [27:0] _T_1219; // @[BTB.scala 293:28]
  wire  _T_1220; // @[BTB.scala 293:72]
  wire [8:0] _GEN_448; // @[BTB.scala 87:42]
  wire [8:0] _T_1227; // @[BTB.scala 87:42]
  wire [15:0] _T_1228; // @[BTB.scala 83:12]
  wire [8:0] _T_1230; // @[BTB.scala 89:44]
  wire [7:0] _T_1235; // @[Cat.scala 30:58]
  wire [8:0] _GEN_449; // @[BTB.scala 87:42]
  wire [8:0] _T_1240; // @[BTB.scala 87:42]
  wire [15:0] _T_1241; // @[BTB.scala 83:12]
  wire [8:0] _T_1243; // @[BTB.scala 89:44]
  wire [7:0] _T_1247; // @[Cat.scala 30:58]
  wire  _T_1222_value; // @[BTB.scala 92:19 BTB.scala 93:15]
  wire  _T_1250; // @[BTB.scala 308:22]
  reg [2:0] _T_1252; // @[BTB.scala 57:26]
  reg [31:0] _RAND_189;
  reg [2:0] _T_1254; // @[BTB.scala 58:24]
  reg [31:0] _RAND_190;
  reg [38:0] _T_1258_0; // @[BTB.scala 59:26]
  reg [63:0] _RAND_191;
  reg [38:0] _T_1258_1; // @[BTB.scala 59:26]
  reg [63:0] _RAND_192;
  reg [38:0] _T_1258_2; // @[BTB.scala 59:26]
  reg [63:0] _RAND_193;
  reg [38:0] _T_1258_3; // @[BTB.scala 59:26]
  reg [63:0] _RAND_194;
  reg [38:0] _T_1258_4; // @[BTB.scala 59:26]
  reg [63:0] _RAND_195;
  reg [38:0] _T_1258_5; // @[BTB.scala 59:26]
  reg [63:0] _RAND_196;
  wire  _T_1267; // @[BTB.scala 314:42]
  wire  _T_1268; // @[BTB.scala 314:42]
  wire  _T_1269; // @[BTB.scala 314:42]
  wire  _T_1270; // @[BTB.scala 314:42]
  wire  _T_1271; // @[BTB.scala 314:42]
  wire  _T_1272; // @[BTB.scala 314:42]
  wire  _T_1273; // @[BTB.scala 314:42]
  wire  _T_1274; // @[BTB.scala 314:42]
  wire  _T_1275; // @[BTB.scala 314:42]
  wire  _T_1276; // @[BTB.scala 314:42]
  wire  _T_1277; // @[BTB.scala 314:42]
  wire  _T_1278; // @[BTB.scala 314:42]
  wire  _T_1279; // @[BTB.scala 314:42]
  wire  _T_1280; // @[BTB.scala 314:42]
  wire  _T_1281; // @[BTB.scala 314:42]
  wire  _T_1282; // @[BTB.scala 314:42]
  wire  _T_1283; // @[BTB.scala 314:42]
  wire  _T_1284; // @[BTB.scala 314:42]
  wire  _T_1285; // @[BTB.scala 314:42]
  wire  _T_1286; // @[BTB.scala 314:42]
  wire  _T_1287; // @[BTB.scala 314:42]
  wire  _T_1288; // @[BTB.scala 314:42]
  wire  _T_1289; // @[BTB.scala 314:42]
  wire  _T_1290; // @[BTB.scala 314:42]
  wire  _T_1291; // @[BTB.scala 314:42]
  wire  _T_1292; // @[BTB.scala 314:42]
  wire  _T_1293; // @[BTB.scala 314:42]
  wire  _T_1294; // @[BTB.scala 314:42]
  wire [6:0] _T_1300; // @[Cat.scala 30:58]
  wire [13:0] _T_1307; // @[Cat.scala 30:58]
  wire [6:0] _T_1313; // @[Cat.scala 30:58]
  wire [27:0] _T_1321; // @[Cat.scala 30:58]
  wire [27:0] _T_1322; // @[BTB.scala 314:26]
  wire  _T_1323; // @[BTB.scala 314:67]
  wire  _T_1324; // @[BTB.scala 55:29]
  wire [38:0] _GEN_399; // @[BTB.scala 316:22]
  wire [38:0] _GEN_400; // @[BTB.scala 316:22]
  wire [38:0] _GEN_401; // @[BTB.scala 316:22]
  wire [38:0] _GEN_402; // @[BTB.scala 316:22]
  wire [38:0] _GEN_403; // @[BTB.scala 316:22]
  wire  _T_1329; // @[BTB.scala 317:24]
  wire  _T_1331; // @[BTB.scala 321:40]
  wire  _T_1332; // @[BTB.scala 44:17]
  wire [2:0] _T_1334; // @[BTB.scala 44:42]
  wire  _T_1335; // @[BTB.scala 45:49]
  wire [2:0] _T_1338; // @[BTB.scala 45:62]
  wire [2:0] _T_1339; // @[BTB.scala 45:22]
  wire  _T_1341; // @[BTB.scala 323:46]
  wire [2:0] _T_1346; // @[BTB.scala 51:20]
  wire  _T_1347; // @[BTB.scala 52:42]
  wire [2:0] _T_1351; // @[BTB.scala 52:50]
  reg [19:0] BTB_state; // @[Register tracking BTB state]
  reg [31:0] _RAND_197;
  reg  BTB_cov [0:1048575]; // @[Coverage map for BTB]
  reg [31:0] _RAND_198;
  wire  BTB_cov_read_data; // @[Coverage map for BTB]
  wire [19:0] BTB_cov_read_addr; // @[Coverage map for BTB]
  wire  BTB_cov_write_data; // @[Coverage map for BTB]
  wire [19:0] BTB_cov_write_addr; // @[Coverage map for BTB]
  wire  BTB_cov_write_mask; // @[Coverage map for BTB]
  wire  BTB_cov_write_en; // @[Coverage map for BTB]
  reg [29:0] BTB_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_199;
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  mux_cond_4;
  wire  mux_cond_5;
  wire  mux_cond_6;
  wire  mux_cond_7;
  wire  mux_cond_8;
  wire  mux_cond_9;
  wire  mux_cond_10;
  wire  mux_cond_11;
  wire  mux_cond_12;
  wire  mux_cond_13;
  wire  mux_cond_14;
  wire  mux_cond_15;
  wire  mux_cond_16;
  wire  mux_cond_17;
  wire  mux_cond_18;
  wire  mux_cond_19;
  wire  mux_cond_20;
  wire  mux_cond_21;
  wire  mux_cond_22;
  wire  mux_cond_23;
  wire  mux_cond_24;
  wire  mux_cond_25;
  wire  mux_cond_26;
  wire  mux_cond_27;
  wire  mux_cond_28;
  wire [5:0] r_resp_bits_taken_shl;
  wire [19:0] r_resp_bits_taken_pad;
  wire [9:0] _T_1252_shl;
  wire [19:0] _T_1252_pad;
  wire [8:0] pageValid_shl;
  wire [19:0] pageValid_pad;
  wire [5:0] r_btb_update_valid_shl;
  wire [19:0] r_btb_update_valid_pad;
  wire [5:0] _T_1254_shl;
  wire [19:0] _T_1254_pad;
  wire [6:0] r_resp_valid_shl;
  wire [19:0] r_resp_valid_pad;
  wire [11:0] r_btb_update_bits_isValid_shl;
  wire [19:0] r_btb_update_bits_isValid_pad;
  wire [7:0] nextPageRepl_shl;
  wire [19:0] nextPageRepl_pad;
  wire [18:0] mux_cond_0_shl;
  wire [19:0] mux_cond_0_pad;
  wire [8:0] mux_cond_1_shl;
  wire [19:0] mux_cond_1_pad;
  wire [15:0] mux_cond_2_shl;
  wire [19:0] mux_cond_2_pad;
  wire [8:0] mux_cond_3_shl;
  wire [19:0] mux_cond_3_pad;
  wire [1:0] mux_cond_4_shl;
  wire [19:0] mux_cond_4_pad;
  wire [11:0] mux_cond_5_shl;
  wire [19:0] mux_cond_5_pad;
  wire [4:0] mux_cond_6_shl;
  wire [19:0] mux_cond_6_pad;
  wire [15:0] mux_cond_7_shl;
  wire [19:0] mux_cond_7_pad;
  wire [19:0] mux_cond_8_shl;
  wire [19:0] mux_cond_8_pad;
  wire [10:0] mux_cond_9_shl;
  wire [19:0] mux_cond_9_pad;
  wire [6:0] mux_cond_10_shl;
  wire [19:0] mux_cond_10_pad;
  wire [4:0] mux_cond_11_shl;
  wire [19:0] mux_cond_11_pad;
  wire [14:0] mux_cond_12_shl;
  wire [19:0] mux_cond_12_pad;
  wire [3:0] mux_cond_13_shl;
  wire [19:0] mux_cond_13_pad;
  wire [17:0] mux_cond_14_shl;
  wire [19:0] mux_cond_14_pad;
  wire [10:0] mux_cond_15_shl;
  wire [19:0] mux_cond_15_pad;
  wire [18:0] mux_cond_16_shl;
  wire [19:0] mux_cond_16_pad;
  wire [17:0] mux_cond_17_shl;
  wire [19:0] mux_cond_17_pad;
  wire [8:0] mux_cond_18_shl;
  wire [19:0] mux_cond_18_pad;
  wire [8:0] mux_cond_19_shl;
  wire [19:0] mux_cond_19_pad;
  wire [3:0] mux_cond_20_shl;
  wire [19:0] mux_cond_20_pad;
  wire [6:0] mux_cond_21_shl;
  wire [19:0] mux_cond_21_pad;
  wire [19:0] mux_cond_22_shl;
  wire [19:0] mux_cond_22_pad;
  wire [10:0] mux_cond_23_shl;
  wire [19:0] mux_cond_23_pad;
  wire [1:0] mux_cond_24_shl;
  wire [19:0] mux_cond_24_pad;
  wire  mux_cond_25_shl;
  wire [19:0] mux_cond_25_pad;
  wire [8:0] mux_cond_26_shl;
  wire [19:0] mux_cond_26_pad;
  wire [2:0] mux_cond_27_shl;
  wire [19:0] mux_cond_27_pad;
  wire [3:0] mux_cond_28_shl;
  wire [19:0] mux_cond_28_pad;
  wire [11:0] cfiType_4_shl;
  wire [19:0] cfiType_4_pad;
  wire [7:0] tgtPages_20_shl;
  wire [19:0] tgtPages_20_pad;
  wire [7:0] tgtPages_17_shl;
  wire [19:0] tgtPages_17_pad;
  wire [7:0] tgtPages_3_shl;
  wire [19:0] tgtPages_3_pad;
  wire [11:0] cfiType_1_shl;
  wire [19:0] cfiType_1_pad;
  wire [7:0] tgtPages_2_shl;
  wire [19:0] tgtPages_2_pad;
  wire [11:0] cfiType_18_shl;
  wire [19:0] cfiType_18_pad;
  wire [7:0] tgtPages_26_shl;
  wire [19:0] tgtPages_26_pad;
  wire [11:0] cfiType_20_shl;
  wire [19:0] cfiType_20_pad;
  wire [11:0] cfiType_22_shl;
  wire [19:0] cfiType_22_pad;
  wire [11:0] cfiType_23_shl;
  wire [19:0] cfiType_23_pad;
  wire [11:0] cfiType_0_shl;
  wire [19:0] cfiType_0_pad;
  wire [7:0] tgtPages_11_shl;
  wire [19:0] tgtPages_11_pad;
  wire [11:0] cfiType_7_shl;
  wire [19:0] cfiType_7_pad;
  wire [11:0] cfiType_19_shl;
  wire [19:0] cfiType_19_pad;
  wire [11:0] cfiType_17_shl;
  wire [19:0] cfiType_17_pad;
  wire [11:0] cfiType_25_shl;
  wire [19:0] cfiType_25_pad;
  wire [11:0] cfiType_3_shl;
  wire [19:0] cfiType_3_pad;
  wire [11:0] cfiType_10_shl;
  wire [19:0] cfiType_10_pad;
  wire [7:0] tgtPages_14_shl;
  wire [19:0] tgtPages_14_pad;
  wire [11:0] cfiType_2_shl;
  wire [19:0] cfiType_2_pad;
  wire [11:0] cfiType_16_shl;
  wire [19:0] cfiType_16_pad;
  wire [7:0] tgtPages_0_shl;
  wire [19:0] tgtPages_0_pad;
  wire [7:0] tgtPages_21_shl;
  wire [19:0] tgtPages_21_pad;
  wire [7:0] tgtPages_5_shl;
  wire [19:0] tgtPages_5_pad;
  wire [7:0] tgtPages_4_shl;
  wire [19:0] tgtPages_4_pad;
  wire [11:0] cfiType_9_shl;
  wire [19:0] cfiType_9_pad;
  wire [7:0] tgtPages_25_shl;
  wire [19:0] tgtPages_25_pad;
  wire [11:0] cfiType_8_shl;
  wire [19:0] cfiType_8_pad;
  wire [7:0] tgtPages_24_shl;
  wire [19:0] tgtPages_24_pad;
  wire [11:0] cfiType_26_shl;
  wire [19:0] cfiType_26_pad;
  wire [7:0] tgtPages_13_shl;
  wire [19:0] tgtPages_13_pad;
  wire [11:0] cfiType_14_shl;
  wire [19:0] cfiType_14_pad;
  wire [11:0] cfiType_11_shl;
  wire [19:0] cfiType_11_pad;
  wire [7:0] tgtPages_16_shl;
  wire [19:0] tgtPages_16_pad;
  wire [11:0] cfiType_15_shl;
  wire [19:0] cfiType_15_pad;
  wire [11:0] cfiType_24_shl;
  wire [19:0] cfiType_24_pad;
  wire [7:0] tgtPages_18_shl;
  wire [19:0] tgtPages_18_pad;
  wire [11:0] cfiType_21_shl;
  wire [19:0] cfiType_21_pad;
  wire [7:0] tgtPages_12_shl;
  wire [19:0] tgtPages_12_pad;
  wire [7:0] tgtPages_10_shl;
  wire [19:0] tgtPages_10_pad;
  wire [7:0] tgtPages_15_shl;
  wire [19:0] tgtPages_15_pad;
  wire [7:0] tgtPages_22_shl;
  wire [19:0] tgtPages_22_pad;
  wire [7:0] tgtPages_19_shl;
  wire [19:0] tgtPages_19_pad;
  wire [11:0] cfiType_13_shl;
  wire [19:0] cfiType_13_pad;
  wire [11:0] cfiType_6_shl;
  wire [19:0] cfiType_6_pad;
  wire [7:0] tgtPages_6_shl;
  wire [19:0] tgtPages_6_pad;
  wire [11:0] cfiType_27_shl;
  wire [19:0] cfiType_27_pad;
  wire [7:0] tgtPages_23_shl;
  wire [19:0] tgtPages_23_pad;
  wire [11:0] cfiType_12_shl;
  wire [19:0] cfiType_12_pad;
  wire [7:0] tgtPages_8_shl;
  wire [19:0] tgtPages_8_pad;
  wire [7:0] tgtPages_1_shl;
  wire [19:0] tgtPages_1_pad;
  wire [7:0] tgtPages_9_shl;
  wire [19:0] tgtPages_9_pad;
  wire [11:0] cfiType_5_shl;
  wire [19:0] cfiType_5_pad;
  wire [7:0] tgtPages_7_shl;
  wire [19:0] tgtPages_7_pad;
  wire [7:0] tgtPages_27_shl;
  wire [19:0] tgtPages_27_pad;
  wire [19:0] BTB_xor31;
  wire [19:0] BTB_xor66;
  wire [19:0] BTB_xor32;
  wire [19:0] BTB_xor15;
  wire [19:0] BTB_xor68;
  wire [19:0] BTB_xor33;
  wire [19:0] BTB_xor70;
  wire [19:0] BTB_xor34;
  wire [19:0] BTB_xor16;
  wire [19:0] BTB_xor7;
  wire [19:0] BTB_xor72;
  wire [19:0] BTB_xor35;
  wire [19:0] BTB_xor74;
  wire [19:0] BTB_xor36;
  wire [19:0] BTB_xor17;
  wire [19:0] BTB_xor76;
  wire [19:0] BTB_xor37;
  wire [19:0] BTB_xor78;
  wire [19:0] BTB_xor38;
  wire [19:0] BTB_xor18;
  wire [19:0] BTB_xor8;
  wire [19:0] BTB_xor3;
  wire [19:0] BTB_xor39;
  wire [19:0] BTB_xor82;
  wire [19:0] BTB_xor40;
  wire [19:0] BTB_xor19;
  wire [19:0] BTB_xor84;
  wire [19:0] BTB_xor41;
  wire [19:0] BTB_xor86;
  wire [19:0] BTB_xor42;
  wire [19:0] BTB_xor20;
  wire [19:0] BTB_xor9;
  wire [19:0] BTB_xor88;
  wire [19:0] BTB_xor43;
  wire [19:0] BTB_xor90;
  wire [19:0] BTB_xor44;
  wire [19:0] BTB_xor21;
  wire [19:0] BTB_xor92;
  wire [19:0] BTB_xor45;
  wire [19:0] BTB_xor94;
  wire [19:0] BTB_xor46;
  wire [19:0] BTB_xor22;
  wire [19:0] BTB_xor10;
  wire [19:0] BTB_xor4;
  wire [19:0] BTB_xor1;
  wire [19:0] BTB_xor47;
  wire [19:0] BTB_xor98;
  wire [19:0] BTB_xor48;
  wire [19:0] BTB_xor23;
  wire [19:0] BTB_xor100;
  wire [19:0] BTB_xor49;
  wire [19:0] BTB_xor102;
  wire [19:0] BTB_xor50;
  wire [19:0] BTB_xor24;
  wire [19:0] BTB_xor11;
  wire [19:0] BTB_xor104;
  wire [19:0] BTB_xor51;
  wire [19:0] BTB_xor106;
  wire [19:0] BTB_xor52;
  wire [19:0] BTB_xor25;
  wire [19:0] BTB_xor108;
  wire [19:0] BTB_xor53;
  wire [19:0] BTB_xor110;
  wire [19:0] BTB_xor54;
  wire [19:0] BTB_xor26;
  wire [19:0] BTB_xor12;
  wire [19:0] BTB_xor5;
  wire [19:0] BTB_xor112;
  wire [19:0] BTB_xor55;
  wire [19:0] BTB_xor114;
  wire [19:0] BTB_xor56;
  wire [19:0] BTB_xor27;
  wire [19:0] BTB_xor116;
  wire [19:0] BTB_xor57;
  wire [19:0] BTB_xor118;
  wire [19:0] BTB_xor58;
  wire [19:0] BTB_xor28;
  wire [19:0] BTB_xor13;
  wire [19:0] BTB_xor120;
  wire [19:0] BTB_xor59;
  wire [19:0] BTB_xor122;
  wire [19:0] BTB_xor60;
  wire [19:0] BTB_xor29;
  wire [19:0] BTB_xor124;
  wire [19:0] BTB_xor61;
  wire [19:0] BTB_xor126;
  wire [19:0] BTB_xor62;
  wire [19:0] BTB_xor30;
  wire [19:0] BTB_xor14;
  wire [19:0] BTB_xor6;
  wire [19:0] BTB_xor2;
  wire [19:0] BTB_xor0;
  assign _T_1161__T_1232_addr = _T_1227 ^ _T_1230;
  assign _T_1161__T_1232_data = _T_1161[_T_1161__T_1232_addr]; // @[BTB.scala 113:26]
  assign _T_1161__T_1245_data = io_bht_update_bits_taken;
  assign _T_1161__T_1245_addr = _T_1240 ^ _T_1243;
  assign _T_1161__T_1245_mask = 1'h1;
  assign _T_1161__T_1245_en = io_bht_update_valid & io_bht_update_bits_branch;
  assign _T_249 = pages_0 == io_req_bits_addr[38:14]; // @[BTB.scala 202:29]
  assign _T_250 = pages_1 == io_req_bits_addr[38:14]; // @[BTB.scala 202:29]
  assign _T_251 = pages_2 == io_req_bits_addr[38:14]; // @[BTB.scala 202:29]
  assign _T_252 = pages_3 == io_req_bits_addr[38:14]; // @[BTB.scala 202:29]
  assign _T_253 = pages_4 == io_req_bits_addr[38:14]; // @[BTB.scala 202:29]
  assign _T_254 = pages_5 == io_req_bits_addr[38:14]; // @[BTB.scala 202:29]
  assign _T_259 = {_T_254,_T_253,_T_252,_T_251,_T_250,_T_249}; // @[Cat.scala 30:58]
  assign pageHit = pageValid & _T_259; // @[BTB.scala 202:15]
  assign _T_261 = idxs_0 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_262 = idxs_1 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_263 = idxs_2 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_264 = idxs_3 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_265 = idxs_4 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_266 = idxs_5 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_267 = idxs_6 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_268 = idxs_7 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_269 = idxs_8 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_270 = idxs_9 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_271 = idxs_10 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_272 = idxs_11 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_273 = idxs_12 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_274 = idxs_13 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_275 = idxs_14 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_276 = idxs_15 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_277 = idxs_16 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_278 = idxs_17 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_279 = idxs_18 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_280 = idxs_19 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_281 = idxs_20 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_282 = idxs_21 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_283 = idxs_22 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_284 = idxs_23 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_285 = idxs_24 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_286 = idxs_25 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_287 = idxs_26 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_288 = idxs_27 == io_req_bits_addr[13:1]; // @[BTB.scala 206:16]
  assign _T_294 = {_T_267,_T_266,_T_265,_T_264,_T_263,_T_262,_T_261}; // @[Cat.scala 30:58]
  assign _T_301 = {_T_274,_T_273,_T_272,_T_271,_T_270,_T_269,_T_268,_T_294}; // @[Cat.scala 30:58]
  assign _T_307 = {_T_281,_T_280,_T_279,_T_278,_T_277,_T_276,_T_275}; // @[Cat.scala 30:58]
  assign _T_315 = {_T_288,_T_287,_T_286,_T_285,_T_284,_T_283,_T_282,_T_307,_T_301}; // @[Cat.scala 30:58]
  assign idxHit = _T_315 & isValid; // @[BTB.scala 206:32]
  assign _T_317 = pages_0 == r_btb_update_bits_pc[38:14]; // @[BTB.scala 202:29]
  assign _T_318 = pages_1 == r_btb_update_bits_pc[38:14]; // @[BTB.scala 202:29]
  assign _T_319 = pages_2 == r_btb_update_bits_pc[38:14]; // @[BTB.scala 202:29]
  assign _T_320 = pages_3 == r_btb_update_bits_pc[38:14]; // @[BTB.scala 202:29]
  assign _T_321 = pages_4 == r_btb_update_bits_pc[38:14]; // @[BTB.scala 202:29]
  assign _T_322 = pages_5 == r_btb_update_bits_pc[38:14]; // @[BTB.scala 202:29]
  assign _T_327 = {_T_322,_T_321,_T_320,_T_319,_T_318,_T_317}; // @[Cat.scala 30:58]
  assign updatePageHit = pageValid & _T_327; // @[BTB.scala 202:15]
  assign updateHit = r_btb_update_bits_prediction_entry < 5'h1c; // @[BTB.scala 220:48]
  assign useUpdatePageHit = updatePageHit != 6'h0; // @[BTB.scala 222:40]
  assign usePageHit = pageHit != 6'h0; // @[BTB.scala 223:28]
  assign doIdxPageRepl = ~useUpdatePageHit; // @[BTB.scala 224:23]
  assign _T_331 = {pageHit[4:0],pageHit[5]}; // @[Cat.scala 30:58]
  assign _T_332 = 8'h1 << nextPageRepl; // @[OneHot.scala 45:35]
  assign _T_333 = usePageHit ? 8'h0 : _T_332; // @[BTB.scala 226:70]
  assign _GEN_432 = {{2'd0}, _T_331}; // @[BTB.scala 226:65]
  assign idxPageRepl = _GEN_432 | _T_333; // @[BTB.scala 226:65]
  assign idxPageUpdateOH = useUpdatePageHit ? {{2'd0}, updatePageHit} : idxPageRepl; // @[BTB.scala 227:28]
  assign _T_336 = idxPageUpdateOH[7:4] != 4'h0; // @[OneHot.scala 28:14]
  assign _T_337 = idxPageUpdateOH[7:4] | idxPageUpdateOH[3:0]; // @[OneHot.scala 28:28]
  assign _T_340 = _T_337[3:2] != 2'h0; // @[OneHot.scala 28:14]
  assign _T_341 = _T_337[3:2] | _T_337[1:0]; // @[OneHot.scala 28:28]
  assign idxPageUpdate = {_T_336,_T_340,_T_341[1]}; // @[Cat.scala 30:58]
  assign idxPageReplEn = doIdxPageRepl ? idxPageRepl : 8'h0; // @[BTB.scala 229:26]
  assign samePage = r_btb_update_bits_pc[38:14] == io_req_bits_addr[38:14]; // @[BTB.scala 231:45]
  assign doTgtPageRepl = ~samePage & ~usePageHit; // @[BTB.scala 232:33]
  assign _T_350 = {idxPageUpdateOH[4:0],idxPageUpdateOH[5]}; // @[Cat.scala 30:58]
  assign tgtPageRepl = samePage ? idxPageUpdateOH : {{2'd0}, _T_350}; // @[BTB.scala 233:24]
  assign _T_351 = usePageHit ? 8'h0 : tgtPageRepl; // @[BTB.scala 234:45]
  assign _GEN_433 = {{2'd0}, pageHit}; // @[BTB.scala 234:40]
  assign _T_352 = _GEN_433 | _T_351; // @[BTB.scala 234:40]
  assign _T_355 = _T_352[7:4] != 4'h0; // @[OneHot.scala 28:14]
  assign _T_356 = _T_352[7:4] | _T_352[3:0]; // @[OneHot.scala 28:28]
  assign _T_359 = _T_356[3:2] != 2'h0; // @[OneHot.scala 28:14]
  assign _T_360 = _T_356[3:2] | _T_356[1:0]; // @[OneHot.scala 28:28]
  assign tgtPageUpdate = {_T_355,_T_359,_T_360[1]}; // @[Cat.scala 30:58]
  assign tgtPageReplEn = doTgtPageRepl ? tgtPageRepl : 8'h0; // @[BTB.scala 235:26]
  assign _T_363 = doIdxPageRepl | doTgtPageRepl; // @[BTB.scala 237:46]
  assign _T_364 = r_btb_update_valid & _T_363; // @[BTB.scala 237:28]
  assign _T_365 = doIdxPageRepl & doTgtPageRepl; // @[BTB.scala 238:30]
  assign _T_366 = _T_365 ? 2'h2 : 2'h1; // @[BTB.scala 239:40]
  assign _GEN_434 = {{1'd0}, _T_366}; // @[BTB.scala 239:29]
  assign _T_368 = nextPageRepl + _GEN_434; // @[BTB.scala 239:29]
  assign _T_369 = _T_368 >= 3'h6; // @[BTB.scala 240:30]
  assign _T_374 = {_T_373, 1'h0}; // @[Replacement.scala 57:31]
  assign _T_378 = {{1'd0}, _T_374[27:1]}; // @[Replacement.scala 61:48]
  assign _T_381 = {1'h1,_T_378[0]}; // @[Cat.scala 30:58]
  assign _T_382 = {1'h1,_T_378[0],4'h8}; // @[Cat.scala 30:58]
  assign _T_384 = _T_382[4:0] < 5'h1c; // @[Replacement.scala 60:70]
  assign _T_385 = _T_374 >> _T_381; // @[Replacement.scala 61:48]
  assign _T_387 = _T_384 & _T_385[0]; // @[Replacement.scala 61:32]
  assign _T_388 = {1'h1,_T_378[0],_T_387}; // @[Cat.scala 30:58]
  assign _T_389 = {1'h1,_T_378[0],_T_387,3'h4}; // @[Cat.scala 30:58]
  assign _T_391 = _T_389[4:0] < 5'h1c; // @[Replacement.scala 60:70]
  assign _T_392 = _T_374 >> _T_388; // @[Replacement.scala 61:48]
  assign _T_394 = _T_391 & _T_392[0]; // @[Replacement.scala 61:32]
  assign _T_395 = {1'h1,_T_378[0],_T_387,_T_394}; // @[Cat.scala 30:58]
  assign _T_396 = {1'h1,_T_378[0],_T_387,_T_394,2'h2}; // @[Cat.scala 30:58]
  assign _T_398 = _T_396[4:0] < 5'h1c; // @[Replacement.scala 60:70]
  assign _T_399 = _T_374 >> _T_395; // @[Replacement.scala 61:48]
  assign _T_401 = _T_398 & _T_399[0]; // @[Replacement.scala 61:32]
  assign _T_402 = {1'h1,_T_378[0],_T_387,_T_394,_T_401}; // @[Cat.scala 30:58]
  assign _T_403 = {1'h1,_T_378[0],_T_387,_T_394,_T_401,1'h1}; // @[Cat.scala 30:58]
  assign _T_405 = _T_403[4:0] < 5'h1c; // @[Replacement.scala 60:70]
  assign _T_406 = _T_374 >> _T_402; // @[Replacement.scala 61:48]
  assign _T_408 = _T_405 & _T_406[0]; // @[Replacement.scala 61:32]
  assign _T_409 = {1'h1,_T_378[0],_T_387,_T_394,_T_401,_T_408}; // @[Cat.scala 30:58]
  assign waddr = updateHit ? r_btb_update_bits_prediction_entry : _T_409[4:0]; // @[BTB.scala 244:18]
  assign _T_419 = r_resp_valid & r_resp_bits_taken; // @[BTB.scala 246:22]
  assign _T_420 = _T_419 | r_btb_update_valid; // @[BTB.scala 246:43]
  assign _T_421 = r_btb_update_valid ? waddr : r_resp_bits_entry; // @[BTB.scala 247:20]
  assign _T_426 = _T_374 | 28'h2; // @[Replacement.scala 50:37]
  assign _T_428 = ~_T_374 | 28'h2; // @[Replacement.scala 50:37]
  assign _T_430 = _T_421[4] ? ~_T_428 : _T_426; // @[Replacement.scala 50:37]
  assign _T_431 = {1'h1,_T_421[4]}; // @[Cat.scala 30:58]
  assign _T_434 = 4'h1 << _T_431; // @[Replacement.scala 50:37]
  assign _GEN_436 = {{24'd0}, _T_434}; // @[Replacement.scala 50:37]
  assign _T_435 = _T_430 | _GEN_436; // @[Replacement.scala 50:37]
  assign _T_437 = ~_T_430 | _GEN_436; // @[Replacement.scala 50:37]
  assign _T_439 = _T_421[3] ? ~_T_437 : _T_435; // @[Replacement.scala 50:37]
  assign _T_440 = {1'h1,_T_421[4],_T_421[3]}; // @[Cat.scala 30:58]
  assign _T_443 = 8'h1 << _T_440; // @[Replacement.scala 50:37]
  assign _GEN_438 = {{20'd0}, _T_443}; // @[Replacement.scala 50:37]
  assign _T_444 = _T_439 | _GEN_438; // @[Replacement.scala 50:37]
  assign _T_446 = ~_T_439 | _GEN_438; // @[Replacement.scala 50:37]
  assign _T_448 = _T_421[2] ? ~_T_446 : _T_444; // @[Replacement.scala 50:37]
  assign _T_449 = {1'h1,_T_421[4],_T_421[3],_T_421[2]}; // @[Cat.scala 30:58]
  assign _T_452 = 16'h1 << _T_449; // @[Replacement.scala 50:37]
  assign _GEN_440 = {{12'd0}, _T_452}; // @[Replacement.scala 50:37]
  assign _T_453 = _T_448 | _GEN_440; // @[Replacement.scala 50:37]
  assign _T_455 = ~_T_448 | _GEN_440; // @[Replacement.scala 50:37]
  assign _T_457 = _T_421[1] ? ~_T_455 : _T_453; // @[Replacement.scala 50:37]
  assign _T_458 = {1'h1,_T_421[4],_T_421[3],_T_421[2],_T_421[1]}; // @[Cat.scala 30:58]
  assign _T_461 = 32'h1 << _T_458; // @[Replacement.scala 50:37]
  assign _GEN_442 = {{4'd0}, _T_457}; // @[Replacement.scala 50:37]
  assign _T_462 = _GEN_442 | _T_461; // @[Replacement.scala 50:37]
  assign _GEN_443 = {{4'd0}, ~_T_457}; // @[Replacement.scala 50:37]
  assign _T_464 = _GEN_443 | _T_461; // @[Replacement.scala 50:37]
  assign _T_466 = _T_421[0] ? ~_T_464 : _T_462; // @[Replacement.scala 50:37]
  assign _T_469 = 32'h1 << waddr; // @[OneHot.scala 45:35]
  assign _T_475 = idxPageUpdate + 3'h1; // @[BTB.scala 254:38]
  assign _GEN_444 = {{4'd0}, isValid}; // @[BTB.scala 257:55]
  assign _T_478 = _GEN_444 | _T_469; // @[BTB.scala 257:55]
  assign _T_480 = _GEN_444 & ~_T_469; // @[BTB.scala 257:71]
  assign _T_481 = r_btb_update_bits_isValid ? _T_478 : _T_480; // @[BTB.scala 257:19]
  assign _T_486 = idxPageUpdate[0] ? tgtPageReplEn : idxPageReplEn; // @[BTB.scala 268:24]
  assign _T_493 = idxPageUpdate[0] ? idxPageReplEn : tgtPageReplEn; // @[BTB.scala 270:24]
  assign _GEN_446 = {{2'd0}, pageValid}; // @[BTB.scala 272:28]
  assign _T_500 = _GEN_446 | tgtPageReplEn; // @[BTB.scala 272:28]
  assign _T_501 = _T_500 | idxPageReplEn; // @[BTB.scala 272:44]
  assign _GEN_338 = r_btb_update_valid ? _T_481 : {{4'd0}, isValid}; // @[BTB.scala 250:29]
  assign _GEN_373 = r_btb_update_valid ? _T_501 : {{2'd0}, pageValid}; // @[BTB.scala 250:29]
  assign _T_502 = {pageHit, 1'h0}; // @[BTB.scala 275:29]
  assign _T_532 = idxHit[0] ? idxPages_0 : 3'h0; // @[Mux.scala 19:72]
  assign _T_533 = idxHit[1] ? idxPages_1 : 3'h0; // @[Mux.scala 19:72]
  assign _T_534 = idxHit[2] ? idxPages_2 : 3'h0; // @[Mux.scala 19:72]
  assign _T_535 = idxHit[3] ? idxPages_3 : 3'h0; // @[Mux.scala 19:72]
  assign _T_536 = idxHit[4] ? idxPages_4 : 3'h0; // @[Mux.scala 19:72]
  assign _T_537 = idxHit[5] ? idxPages_5 : 3'h0; // @[Mux.scala 19:72]
  assign _T_538 = idxHit[6] ? idxPages_6 : 3'h0; // @[Mux.scala 19:72]
  assign _T_539 = idxHit[7] ? idxPages_7 : 3'h0; // @[Mux.scala 19:72]
  assign _T_540 = idxHit[8] ? idxPages_8 : 3'h0; // @[Mux.scala 19:72]
  assign _T_541 = idxHit[9] ? idxPages_9 : 3'h0; // @[Mux.scala 19:72]
  assign _T_542 = idxHit[10] ? idxPages_10 : 3'h0; // @[Mux.scala 19:72]
  assign _T_543 = idxHit[11] ? idxPages_11 : 3'h0; // @[Mux.scala 19:72]
  assign _T_544 = idxHit[12] ? idxPages_12 : 3'h0; // @[Mux.scala 19:72]
  assign _T_545 = idxHit[13] ? idxPages_13 : 3'h0; // @[Mux.scala 19:72]
  assign _T_546 = idxHit[14] ? idxPages_14 : 3'h0; // @[Mux.scala 19:72]
  assign _T_547 = idxHit[15] ? idxPages_15 : 3'h0; // @[Mux.scala 19:72]
  assign _T_548 = idxHit[16] ? idxPages_16 : 3'h0; // @[Mux.scala 19:72]
  assign _T_549 = idxHit[17] ? idxPages_17 : 3'h0; // @[Mux.scala 19:72]
  assign _T_550 = idxHit[18] ? idxPages_18 : 3'h0; // @[Mux.scala 19:72]
  assign _T_551 = idxHit[19] ? idxPages_19 : 3'h0; // @[Mux.scala 19:72]
  assign _T_552 = idxHit[20] ? idxPages_20 : 3'h0; // @[Mux.scala 19:72]
  assign _T_553 = idxHit[21] ? idxPages_21 : 3'h0; // @[Mux.scala 19:72]
  assign _T_554 = idxHit[22] ? idxPages_22 : 3'h0; // @[Mux.scala 19:72]
  assign _T_555 = idxHit[23] ? idxPages_23 : 3'h0; // @[Mux.scala 19:72]
  assign _T_556 = idxHit[24] ? idxPages_24 : 3'h0; // @[Mux.scala 19:72]
  assign _T_557 = idxHit[25] ? idxPages_25 : 3'h0; // @[Mux.scala 19:72]
  assign _T_558 = idxHit[26] ? idxPages_26 : 3'h0; // @[Mux.scala 19:72]
  assign _T_559 = idxHit[27] ? idxPages_27 : 3'h0; // @[Mux.scala 19:72]
  assign _T_560 = _T_532 | _T_533; // @[Mux.scala 19:72]
  assign _T_561 = _T_560 | _T_534; // @[Mux.scala 19:72]
  assign _T_562 = _T_561 | _T_535; // @[Mux.scala 19:72]
  assign _T_563 = _T_562 | _T_536; // @[Mux.scala 19:72]
  assign _T_564 = _T_563 | _T_537; // @[Mux.scala 19:72]
  assign _T_565 = _T_564 | _T_538; // @[Mux.scala 19:72]
  assign _T_566 = _T_565 | _T_539; // @[Mux.scala 19:72]
  assign _T_567 = _T_566 | _T_540; // @[Mux.scala 19:72]
  assign _T_568 = _T_567 | _T_541; // @[Mux.scala 19:72]
  assign _T_569 = _T_568 | _T_542; // @[Mux.scala 19:72]
  assign _T_570 = _T_569 | _T_543; // @[Mux.scala 19:72]
  assign _T_571 = _T_570 | _T_544; // @[Mux.scala 19:72]
  assign _T_572 = _T_571 | _T_545; // @[Mux.scala 19:72]
  assign _T_573 = _T_572 | _T_546; // @[Mux.scala 19:72]
  assign _T_574 = _T_573 | _T_547; // @[Mux.scala 19:72]
  assign _T_575 = _T_574 | _T_548; // @[Mux.scala 19:72]
  assign _T_576 = _T_575 | _T_549; // @[Mux.scala 19:72]
  assign _T_577 = _T_576 | _T_550; // @[Mux.scala 19:72]
  assign _T_578 = _T_577 | _T_551; // @[Mux.scala 19:72]
  assign _T_579 = _T_578 | _T_552; // @[Mux.scala 19:72]
  assign _T_580 = _T_579 | _T_553; // @[Mux.scala 19:72]
  assign _T_581 = _T_580 | _T_554; // @[Mux.scala 19:72]
  assign _T_582 = _T_581 | _T_555; // @[Mux.scala 19:72]
  assign _T_583 = _T_582 | _T_556; // @[Mux.scala 19:72]
  assign _T_584 = _T_583 | _T_557; // @[Mux.scala 19:72]
  assign _T_585 = _T_584 | _T_558; // @[Mux.scala 19:72]
  assign _T_586 = _T_585 | _T_559; // @[Mux.scala 19:72]
  assign _T_589 = _T_502 >> _T_586; // @[BTB.scala 275:34]
  assign _T_620 = idxHit[0] ? tgtPages_0 : 3'h0; // @[Mux.scala 19:72]
  assign _T_621 = idxHit[1] ? tgtPages_1 : 3'h0; // @[Mux.scala 19:72]
  assign _T_622 = idxHit[2] ? tgtPages_2 : 3'h0; // @[Mux.scala 19:72]
  assign _T_623 = idxHit[3] ? tgtPages_3 : 3'h0; // @[Mux.scala 19:72]
  assign _T_624 = idxHit[4] ? tgtPages_4 : 3'h0; // @[Mux.scala 19:72]
  assign _T_625 = idxHit[5] ? tgtPages_5 : 3'h0; // @[Mux.scala 19:72]
  assign _T_626 = idxHit[6] ? tgtPages_6 : 3'h0; // @[Mux.scala 19:72]
  assign _T_627 = idxHit[7] ? tgtPages_7 : 3'h0; // @[Mux.scala 19:72]
  assign _T_628 = idxHit[8] ? tgtPages_8 : 3'h0; // @[Mux.scala 19:72]
  assign _T_629 = idxHit[9] ? tgtPages_9 : 3'h0; // @[Mux.scala 19:72]
  assign _T_630 = idxHit[10] ? tgtPages_10 : 3'h0; // @[Mux.scala 19:72]
  assign _T_631 = idxHit[11] ? tgtPages_11 : 3'h0; // @[Mux.scala 19:72]
  assign _T_632 = idxHit[12] ? tgtPages_12 : 3'h0; // @[Mux.scala 19:72]
  assign _T_633 = idxHit[13] ? tgtPages_13 : 3'h0; // @[Mux.scala 19:72]
  assign _T_634 = idxHit[14] ? tgtPages_14 : 3'h0; // @[Mux.scala 19:72]
  assign _T_635 = idxHit[15] ? tgtPages_15 : 3'h0; // @[Mux.scala 19:72]
  assign _T_636 = idxHit[16] ? tgtPages_16 : 3'h0; // @[Mux.scala 19:72]
  assign _T_637 = idxHit[17] ? tgtPages_17 : 3'h0; // @[Mux.scala 19:72]
  assign _T_638 = idxHit[18] ? tgtPages_18 : 3'h0; // @[Mux.scala 19:72]
  assign _T_639 = idxHit[19] ? tgtPages_19 : 3'h0; // @[Mux.scala 19:72]
  assign _T_640 = idxHit[20] ? tgtPages_20 : 3'h0; // @[Mux.scala 19:72]
  assign _T_641 = idxHit[21] ? tgtPages_21 : 3'h0; // @[Mux.scala 19:72]
  assign _T_642 = idxHit[22] ? tgtPages_22 : 3'h0; // @[Mux.scala 19:72]
  assign _T_643 = idxHit[23] ? tgtPages_23 : 3'h0; // @[Mux.scala 19:72]
  assign _T_644 = idxHit[24] ? tgtPages_24 : 3'h0; // @[Mux.scala 19:72]
  assign _T_645 = idxHit[25] ? tgtPages_25 : 3'h0; // @[Mux.scala 19:72]
  assign _T_646 = idxHit[26] ? tgtPages_26 : 3'h0; // @[Mux.scala 19:72]
  assign _T_647 = idxHit[27] ? tgtPages_27 : 3'h0; // @[Mux.scala 19:72]
  assign _T_648 = _T_620 | _T_621; // @[Mux.scala 19:72]
  assign _T_649 = _T_648 | _T_622; // @[Mux.scala 19:72]
  assign _T_650 = _T_649 | _T_623; // @[Mux.scala 19:72]
  assign _T_651 = _T_650 | _T_624; // @[Mux.scala 19:72]
  assign _T_652 = _T_651 | _T_625; // @[Mux.scala 19:72]
  assign _T_653 = _T_652 | _T_626; // @[Mux.scala 19:72]
  assign _T_654 = _T_653 | _T_627; // @[Mux.scala 19:72]
  assign _T_655 = _T_654 | _T_628; // @[Mux.scala 19:72]
  assign _T_656 = _T_655 | _T_629; // @[Mux.scala 19:72]
  assign _T_657 = _T_656 | _T_630; // @[Mux.scala 19:72]
  assign _T_658 = _T_657 | _T_631; // @[Mux.scala 19:72]
  assign _T_659 = _T_658 | _T_632; // @[Mux.scala 19:72]
  assign _T_660 = _T_659 | _T_633; // @[Mux.scala 19:72]
  assign _T_661 = _T_660 | _T_634; // @[Mux.scala 19:72]
  assign _T_662 = _T_661 | _T_635; // @[Mux.scala 19:72]
  assign _T_663 = _T_662 | _T_636; // @[Mux.scala 19:72]
  assign _T_664 = _T_663 | _T_637; // @[Mux.scala 19:72]
  assign _T_665 = _T_664 | _T_638; // @[Mux.scala 19:72]
  assign _T_666 = _T_665 | _T_639; // @[Mux.scala 19:72]
  assign _T_667 = _T_666 | _T_640; // @[Mux.scala 19:72]
  assign _T_668 = _T_667 | _T_641; // @[Mux.scala 19:72]
  assign _T_669 = _T_668 | _T_642; // @[Mux.scala 19:72]
  assign _T_670 = _T_669 | _T_643; // @[Mux.scala 19:72]
  assign _T_671 = _T_670 | _T_644; // @[Mux.scala 19:72]
  assign _T_672 = _T_671 | _T_645; // @[Mux.scala 19:72]
  assign _T_673 = _T_672 | _T_646; // @[Mux.scala 19:72]
  assign _T_674 = _T_673 | _T_647; // @[Mux.scala 19:72]
  assign _T_707 = idxHit[0] ? tgts_0 : 13'h0; // @[Mux.scala 19:72]
  assign _T_708 = idxHit[1] ? tgts_1 : 13'h0; // @[Mux.scala 19:72]
  assign _T_709 = idxHit[2] ? tgts_2 : 13'h0; // @[Mux.scala 19:72]
  assign _T_710 = idxHit[3] ? tgts_3 : 13'h0; // @[Mux.scala 19:72]
  assign _T_711 = idxHit[4] ? tgts_4 : 13'h0; // @[Mux.scala 19:72]
  assign _T_712 = idxHit[5] ? tgts_5 : 13'h0; // @[Mux.scala 19:72]
  assign _T_713 = idxHit[6] ? tgts_6 : 13'h0; // @[Mux.scala 19:72]
  assign _T_714 = idxHit[7] ? tgts_7 : 13'h0; // @[Mux.scala 19:72]
  assign _T_715 = idxHit[8] ? tgts_8 : 13'h0; // @[Mux.scala 19:72]
  assign _T_716 = idxHit[9] ? tgts_9 : 13'h0; // @[Mux.scala 19:72]
  assign _T_717 = idxHit[10] ? tgts_10 : 13'h0; // @[Mux.scala 19:72]
  assign _T_718 = idxHit[11] ? tgts_11 : 13'h0; // @[Mux.scala 19:72]
  assign _T_719 = idxHit[12] ? tgts_12 : 13'h0; // @[Mux.scala 19:72]
  assign _T_720 = idxHit[13] ? tgts_13 : 13'h0; // @[Mux.scala 19:72]
  assign _T_721 = idxHit[14] ? tgts_14 : 13'h0; // @[Mux.scala 19:72]
  assign _T_722 = idxHit[15] ? tgts_15 : 13'h0; // @[Mux.scala 19:72]
  assign _T_723 = idxHit[16] ? tgts_16 : 13'h0; // @[Mux.scala 19:72]
  assign _T_724 = idxHit[17] ? tgts_17 : 13'h0; // @[Mux.scala 19:72]
  assign _T_725 = idxHit[18] ? tgts_18 : 13'h0; // @[Mux.scala 19:72]
  assign _T_726 = idxHit[19] ? tgts_19 : 13'h0; // @[Mux.scala 19:72]
  assign _T_727 = idxHit[20] ? tgts_20 : 13'h0; // @[Mux.scala 19:72]
  assign _T_728 = idxHit[21] ? tgts_21 : 13'h0; // @[Mux.scala 19:72]
  assign _T_729 = idxHit[22] ? tgts_22 : 13'h0; // @[Mux.scala 19:72]
  assign _T_730 = idxHit[23] ? tgts_23 : 13'h0; // @[Mux.scala 19:72]
  assign _T_731 = idxHit[24] ? tgts_24 : 13'h0; // @[Mux.scala 19:72]
  assign _T_732 = idxHit[25] ? tgts_25 : 13'h0; // @[Mux.scala 19:72]
  assign _T_733 = idxHit[26] ? tgts_26 : 13'h0; // @[Mux.scala 19:72]
  assign _T_734 = idxHit[27] ? tgts_27 : 13'h0; // @[Mux.scala 19:72]
  assign _T_735 = _T_707 | _T_708; // @[Mux.scala 19:72]
  assign _T_736 = _T_735 | _T_709; // @[Mux.scala 19:72]
  assign _T_737 = _T_736 | _T_710; // @[Mux.scala 19:72]
  assign _T_738 = _T_737 | _T_711; // @[Mux.scala 19:72]
  assign _T_739 = _T_738 | _T_712; // @[Mux.scala 19:72]
  assign _T_740 = _T_739 | _T_713; // @[Mux.scala 19:72]
  assign _T_741 = _T_740 | _T_714; // @[Mux.scala 19:72]
  assign _T_742 = _T_741 | _T_715; // @[Mux.scala 19:72]
  assign _T_743 = _T_742 | _T_716; // @[Mux.scala 19:72]
  assign _T_744 = _T_743 | _T_717; // @[Mux.scala 19:72]
  assign _T_745 = _T_744 | _T_718; // @[Mux.scala 19:72]
  assign _T_746 = _T_745 | _T_719; // @[Mux.scala 19:72]
  assign _T_747 = _T_746 | _T_720; // @[Mux.scala 19:72]
  assign _T_748 = _T_747 | _T_721; // @[Mux.scala 19:72]
  assign _T_749 = _T_748 | _T_722; // @[Mux.scala 19:72]
  assign _T_750 = _T_749 | _T_723; // @[Mux.scala 19:72]
  assign _T_751 = _T_750 | _T_724; // @[Mux.scala 19:72]
  assign _T_752 = _T_751 | _T_725; // @[Mux.scala 19:72]
  assign _T_753 = _T_752 | _T_726; // @[Mux.scala 19:72]
  assign _T_754 = _T_753 | _T_727; // @[Mux.scala 19:72]
  assign _T_755 = _T_754 | _T_728; // @[Mux.scala 19:72]
  assign _T_756 = _T_755 | _T_729; // @[Mux.scala 19:72]
  assign _T_757 = _T_756 | _T_730; // @[Mux.scala 19:72]
  assign _T_758 = _T_757 | _T_731; // @[Mux.scala 19:72]
  assign _T_759 = _T_758 | _T_732; // @[Mux.scala 19:72]
  assign _T_760 = _T_759 | _T_733; // @[Mux.scala 19:72]
  assign _T_761 = _T_760 | _T_734; // @[Mux.scala 19:72]
  assign _T_764 = {_T_761, 1'h0}; // @[BTB.scala 277:82]
  assign _GEN_375 = 3'h1 == _T_674 ? pages_1 : pages_0; // @[Cat.scala 30:58]
  assign _GEN_376 = 3'h2 == _T_674 ? pages_2 : _GEN_375; // @[Cat.scala 30:58]
  assign _GEN_377 = 3'h3 == _T_674 ? pages_3 : _GEN_376; // @[Cat.scala 30:58]
  assign _GEN_378 = 3'h4 == _T_674 ? pages_4 : _GEN_377; // @[Cat.scala 30:58]
  assign _GEN_379 = 3'h5 == _T_674 ? pages_5 : _GEN_378; // @[Cat.scala 30:58]
  assign _T_765 = {_GEN_379,_T_764}; // @[Cat.scala 30:58]
  assign _T_768 = idxHit[27:16] != 12'h0; // @[OneHot.scala 28:14]
  assign _GEN_447 = {{4'd0}, idxHit[27:16]}; // @[OneHot.scala 28:28]
  assign _T_769 = _GEN_447 | idxHit[15:0]; // @[OneHot.scala 28:28]
  assign _T_772 = _T_769[15:8] != 8'h0; // @[OneHot.scala 28:14]
  assign _T_773 = _T_769[15:8] | _T_769[7:0]; // @[OneHot.scala 28:28]
  assign _T_776 = _T_773[7:4] != 4'h0; // @[OneHot.scala 28:14]
  assign _T_777 = _T_773[7:4] | _T_773[3:0]; // @[OneHot.scala 28:28]
  assign _T_780 = _T_777[3:2] != 2'h0; // @[OneHot.scala 28:14]
  assign _T_781 = _T_777[3:2] | _T_777[1:0]; // @[OneHot.scala 28:28]
  assign _T_785 = {_T_772,_T_776,_T_780,_T_781[1]}; // @[Cat.scala 30:58]
  assign _T_816 = idxHit[0] & brIdx_0; // @[Mux.scala 19:72]
  assign _T_817 = idxHit[1] & brIdx_1; // @[Mux.scala 19:72]
  assign _T_818 = idxHit[2] & brIdx_2; // @[Mux.scala 19:72]
  assign _T_819 = idxHit[3] & brIdx_3; // @[Mux.scala 19:72]
  assign _T_820 = idxHit[4] & brIdx_4; // @[Mux.scala 19:72]
  assign _T_821 = idxHit[5] & brIdx_5; // @[Mux.scala 19:72]
  assign _T_822 = idxHit[6] & brIdx_6; // @[Mux.scala 19:72]
  assign _T_823 = idxHit[7] & brIdx_7; // @[Mux.scala 19:72]
  assign _T_824 = idxHit[8] & brIdx_8; // @[Mux.scala 19:72]
  assign _T_825 = idxHit[9] & brIdx_9; // @[Mux.scala 19:72]
  assign _T_826 = idxHit[10] & brIdx_10; // @[Mux.scala 19:72]
  assign _T_827 = idxHit[11] & brIdx_11; // @[Mux.scala 19:72]
  assign _T_828 = idxHit[12] & brIdx_12; // @[Mux.scala 19:72]
  assign _T_829 = idxHit[13] & brIdx_13; // @[Mux.scala 19:72]
  assign _T_830 = idxHit[14] & brIdx_14; // @[Mux.scala 19:72]
  assign _T_831 = idxHit[15] & brIdx_15; // @[Mux.scala 19:72]
  assign _T_832 = idxHit[16] & brIdx_16; // @[Mux.scala 19:72]
  assign _T_833 = idxHit[17] & brIdx_17; // @[Mux.scala 19:72]
  assign _T_834 = idxHit[18] & brIdx_18; // @[Mux.scala 19:72]
  assign _T_835 = idxHit[19] & brIdx_19; // @[Mux.scala 19:72]
  assign _T_836 = idxHit[20] & brIdx_20; // @[Mux.scala 19:72]
  assign _T_837 = idxHit[21] & brIdx_21; // @[Mux.scala 19:72]
  assign _T_838 = idxHit[22] & brIdx_22; // @[Mux.scala 19:72]
  assign _T_839 = idxHit[23] & brIdx_23; // @[Mux.scala 19:72]
  assign _T_840 = idxHit[24] & brIdx_24; // @[Mux.scala 19:72]
  assign _T_841 = idxHit[25] & brIdx_25; // @[Mux.scala 19:72]
  assign _T_842 = idxHit[26] & brIdx_26; // @[Mux.scala 19:72]
  assign _T_843 = idxHit[27] & brIdx_27; // @[Mux.scala 19:72]
  assign _T_844 = _T_816 | _T_817; // @[Mux.scala 19:72]
  assign _T_845 = _T_844 | _T_818; // @[Mux.scala 19:72]
  assign _T_846 = _T_845 | _T_819; // @[Mux.scala 19:72]
  assign _T_847 = _T_846 | _T_820; // @[Mux.scala 19:72]
  assign _T_848 = _T_847 | _T_821; // @[Mux.scala 19:72]
  assign _T_849 = _T_848 | _T_822; // @[Mux.scala 19:72]
  assign _T_850 = _T_849 | _T_823; // @[Mux.scala 19:72]
  assign _T_851 = _T_850 | _T_824; // @[Mux.scala 19:72]
  assign _T_852 = _T_851 | _T_825; // @[Mux.scala 19:72]
  assign _T_853 = _T_852 | _T_826; // @[Mux.scala 19:72]
  assign _T_854 = _T_853 | _T_827; // @[Mux.scala 19:72]
  assign _T_855 = _T_854 | _T_828; // @[Mux.scala 19:72]
  assign _T_856 = _T_855 | _T_829; // @[Mux.scala 19:72]
  assign _T_857 = _T_856 | _T_830; // @[Mux.scala 19:72]
  assign _T_858 = _T_857 | _T_831; // @[Mux.scala 19:72]
  assign _T_859 = _T_858 | _T_832; // @[Mux.scala 19:72]
  assign _T_860 = _T_859 | _T_833; // @[Mux.scala 19:72]
  assign _T_861 = _T_860 | _T_834; // @[Mux.scala 19:72]
  assign _T_862 = _T_861 | _T_835; // @[Mux.scala 19:72]
  assign _T_863 = _T_862 | _T_836; // @[Mux.scala 19:72]
  assign _T_864 = _T_863 | _T_837; // @[Mux.scala 19:72]
  assign _T_865 = _T_864 | _T_838; // @[Mux.scala 19:72]
  assign _T_866 = _T_865 | _T_839; // @[Mux.scala 19:72]
  assign _T_867 = _T_866 | _T_840; // @[Mux.scala 19:72]
  assign _T_868 = _T_867 | _T_841; // @[Mux.scala 19:72]
  assign _T_869 = _T_868 | _T_842; // @[Mux.scala 19:72]
  assign _T_977 = idxHit[1] | idxHit[2]; // @[Misc.scala 187:16]
  assign _T_979 = idxHit[1] & idxHit[2]; // @[Misc.scala 187:61]
  assign _T_981 = idxHit[0] | _T_977; // @[Misc.scala 187:16]
  assign _T_983 = idxHit[0] & _T_977; // @[Misc.scala 187:61]
  assign _T_984 = _T_979 | _T_983; // @[Misc.scala 187:49]
  assign _T_991 = idxHit[3] | idxHit[4]; // @[Misc.scala 187:16]
  assign _T_993 = idxHit[3] & idxHit[4]; // @[Misc.scala 187:61]
  assign _T_1000 = idxHit[5] | idxHit[6]; // @[Misc.scala 187:16]
  assign _T_1002 = idxHit[5] & idxHit[6]; // @[Misc.scala 187:61]
  assign _T_1004 = _T_991 | _T_1000; // @[Misc.scala 187:16]
  assign _T_1005 = _T_993 | _T_1002; // @[Misc.scala 187:37]
  assign _T_1006 = _T_991 & _T_1000; // @[Misc.scala 187:61]
  assign _T_1007 = _T_1005 | _T_1006; // @[Misc.scala 187:49]
  assign _T_1008 = _T_981 | _T_1004; // @[Misc.scala 187:16]
  assign _T_1009 = _T_984 | _T_1007; // @[Misc.scala 187:37]
  assign _T_1010 = _T_981 & _T_1004; // @[Misc.scala 187:61]
  assign _T_1011 = _T_1009 | _T_1010; // @[Misc.scala 187:49]
  assign _T_1021 = idxHit[8] | idxHit[9]; // @[Misc.scala 187:16]
  assign _T_1023 = idxHit[8] & idxHit[9]; // @[Misc.scala 187:61]
  assign _T_1025 = idxHit[7] | _T_1021; // @[Misc.scala 187:16]
  assign _T_1027 = idxHit[7] & _T_1021; // @[Misc.scala 187:61]
  assign _T_1028 = _T_1023 | _T_1027; // @[Misc.scala 187:49]
  assign _T_1035 = idxHit[10] | idxHit[11]; // @[Misc.scala 187:16]
  assign _T_1037 = idxHit[10] & idxHit[11]; // @[Misc.scala 187:61]
  assign _T_1044 = idxHit[12] | idxHit[13]; // @[Misc.scala 187:16]
  assign _T_1046 = idxHit[12] & idxHit[13]; // @[Misc.scala 187:61]
  assign _T_1048 = _T_1035 | _T_1044; // @[Misc.scala 187:16]
  assign _T_1049 = _T_1037 | _T_1046; // @[Misc.scala 187:37]
  assign _T_1050 = _T_1035 & _T_1044; // @[Misc.scala 187:61]
  assign _T_1051 = _T_1049 | _T_1050; // @[Misc.scala 187:49]
  assign _T_1052 = _T_1025 | _T_1048; // @[Misc.scala 187:16]
  assign _T_1053 = _T_1028 | _T_1051; // @[Misc.scala 187:37]
  assign _T_1054 = _T_1025 & _T_1048; // @[Misc.scala 187:61]
  assign _T_1055 = _T_1053 | _T_1054; // @[Misc.scala 187:49]
  assign _T_1056 = _T_1008 | _T_1052; // @[Misc.scala 187:16]
  assign _T_1057 = _T_1011 | _T_1055; // @[Misc.scala 187:37]
  assign _T_1058 = _T_1008 & _T_1052; // @[Misc.scala 187:61]
  assign _T_1059 = _T_1057 | _T_1058; // @[Misc.scala 187:49]
  assign _T_1070 = idxHit[15] | idxHit[16]; // @[Misc.scala 187:16]
  assign _T_1072 = idxHit[15] & idxHit[16]; // @[Misc.scala 187:61]
  assign _T_1074 = idxHit[14] | _T_1070; // @[Misc.scala 187:16]
  assign _T_1076 = idxHit[14] & _T_1070; // @[Misc.scala 187:61]
  assign _T_1077 = _T_1072 | _T_1076; // @[Misc.scala 187:49]
  assign _T_1084 = idxHit[17] | idxHit[18]; // @[Misc.scala 187:16]
  assign _T_1086 = idxHit[17] & idxHit[18]; // @[Misc.scala 187:61]
  assign _T_1093 = idxHit[19] | idxHit[20]; // @[Misc.scala 187:16]
  assign _T_1095 = idxHit[19] & idxHit[20]; // @[Misc.scala 187:61]
  assign _T_1097 = _T_1084 | _T_1093; // @[Misc.scala 187:16]
  assign _T_1098 = _T_1086 | _T_1095; // @[Misc.scala 187:37]
  assign _T_1099 = _T_1084 & _T_1093; // @[Misc.scala 187:61]
  assign _T_1100 = _T_1098 | _T_1099; // @[Misc.scala 187:49]
  assign _T_1101 = _T_1074 | _T_1097; // @[Misc.scala 187:16]
  assign _T_1102 = _T_1077 | _T_1100; // @[Misc.scala 187:37]
  assign _T_1103 = _T_1074 & _T_1097; // @[Misc.scala 187:61]
  assign _T_1104 = _T_1102 | _T_1103; // @[Misc.scala 187:49]
  assign _T_1114 = idxHit[22] | idxHit[23]; // @[Misc.scala 187:16]
  assign _T_1116 = idxHit[22] & idxHit[23]; // @[Misc.scala 187:61]
  assign _T_1118 = idxHit[21] | _T_1114; // @[Misc.scala 187:16]
  assign _T_1120 = idxHit[21] & _T_1114; // @[Misc.scala 187:61]
  assign _T_1121 = _T_1116 | _T_1120; // @[Misc.scala 187:49]
  assign _T_1128 = idxHit[24] | idxHit[25]; // @[Misc.scala 187:16]
  assign _T_1130 = idxHit[24] & idxHit[25]; // @[Misc.scala 187:61]
  assign _T_1137 = idxHit[26] | idxHit[27]; // @[Misc.scala 187:16]
  assign _T_1139 = idxHit[26] & idxHit[27]; // @[Misc.scala 187:61]
  assign _T_1141 = _T_1128 | _T_1137; // @[Misc.scala 187:16]
  assign _T_1142 = _T_1130 | _T_1139; // @[Misc.scala 187:37]
  assign _T_1143 = _T_1128 & _T_1137; // @[Misc.scala 187:61]
  assign _T_1144 = _T_1142 | _T_1143; // @[Misc.scala 187:49]
  assign _T_1145 = _T_1118 | _T_1141; // @[Misc.scala 187:16]
  assign _T_1146 = _T_1121 | _T_1144; // @[Misc.scala 187:37]
  assign _T_1147 = _T_1118 & _T_1141; // @[Misc.scala 187:61]
  assign _T_1148 = _T_1146 | _T_1147; // @[Misc.scala 187:49]
  assign _T_1149 = _T_1101 | _T_1145; // @[Misc.scala 187:16]
  assign _T_1150 = _T_1104 | _T_1148; // @[Misc.scala 187:37]
  assign _T_1151 = _T_1101 & _T_1145; // @[Misc.scala 187:61]
  assign _T_1152 = _T_1150 | _T_1151; // @[Misc.scala 187:49]
  assign _T_1154 = _T_1059 | _T_1152; // @[Misc.scala 187:37]
  assign _T_1155 = _T_1056 & _T_1149; // @[Misc.scala 187:61]
  assign _T_1156 = _T_1154 | _T_1155; // @[Misc.scala 187:49]
  assign _T_1158 = isValid & ~idxHit; // @[BTB.scala 285:24]
  assign _GEN_380 = _T_1156 ? {{4'd0}, _T_1158} : _GEN_338; // @[BTB.scala 284:37]
  assign _GEN_381 = io_flush ? 32'h0 : _GEN_380; // @[BTB.scala 287:19]
  assign _T_1164 = cfiType_0 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1165 = cfiType_1 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1166 = cfiType_2 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1167 = cfiType_3 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1168 = cfiType_4 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1169 = cfiType_5 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1170 = cfiType_6 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1171 = cfiType_7 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1172 = cfiType_8 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1173 = cfiType_9 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1174 = cfiType_10 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1175 = cfiType_11 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1176 = cfiType_12 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1177 = cfiType_13 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1178 = cfiType_14 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1179 = cfiType_15 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1180 = cfiType_16 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1181 = cfiType_17 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1182 = cfiType_18 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1183 = cfiType_19 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1184 = cfiType_20 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1185 = cfiType_21 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1186 = cfiType_22 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1187 = cfiType_23 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1188 = cfiType_24 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1189 = cfiType_25 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1190 = cfiType_26 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1191 = cfiType_27 == 2'h0; // @[BTB.scala 293:44]
  assign _T_1197 = {_T_1170,_T_1169,_T_1168,_T_1167,_T_1166,_T_1165,_T_1164}; // @[Cat.scala 30:58]
  assign _T_1204 = {_T_1177,_T_1176,_T_1175,_T_1174,_T_1173,_T_1172,_T_1171,_T_1197}; // @[Cat.scala 30:58]
  assign _T_1210 = {_T_1184,_T_1183,_T_1182,_T_1181,_T_1180,_T_1179,_T_1178}; // @[Cat.scala 30:58]
  assign _T_1218 = {_T_1191,_T_1190,_T_1189,_T_1188,_T_1187,_T_1186,_T_1185,_T_1210,_T_1204}; // @[Cat.scala 30:58]
  assign _T_1219 = idxHit & _T_1218; // @[BTB.scala 293:28]
  assign _T_1220 = _T_1219 != 28'h0; // @[BTB.scala 293:72]
  assign _GEN_448 = {{7'd0}, io_req_bits_addr[12:11]}; // @[BTB.scala 87:42]
  assign _T_1227 = io_req_bits_addr[10:2] ^ _GEN_448; // @[BTB.scala 87:42]
  assign _T_1228 = 8'hdd * _T_1163; // @[BTB.scala 83:12]
  assign _T_1230 = {_T_1228[7:5], 6'h0}; // @[BTB.scala 89:44]
  assign _T_1235 = {io_bht_advance_bits_bht_value,_T_1163[7:1]}; // @[Cat.scala 30:58]
  assign _GEN_449 = {{7'd0}, io_bht_update_bits_pc[12:11]}; // @[BTB.scala 87:42]
  assign _T_1240 = io_bht_update_bits_pc[10:2] ^ _GEN_449; // @[BTB.scala 87:42]
  assign _T_1241 = 8'hdd * io_bht_update_bits_prediction_history; // @[BTB.scala 83:12]
  assign _T_1243 = {_T_1241[7:5], 6'h0}; // @[BTB.scala 89:44]
  assign _T_1247 = {io_bht_update_bits_taken,io_bht_update_bits_prediction_history[7:1]}; // @[Cat.scala 30:58]
  assign _T_1222_value = _T_1161__T_1232_data; // @[BTB.scala 92:19 BTB.scala 93:15]
  assign _T_1250 = ~_T_1222_value & _T_1220; // @[BTB.scala 308:22]
  assign _T_1267 = cfiType_0 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1268 = cfiType_1 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1269 = cfiType_2 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1270 = cfiType_3 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1271 = cfiType_4 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1272 = cfiType_5 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1273 = cfiType_6 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1274 = cfiType_7 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1275 = cfiType_8 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1276 = cfiType_9 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1277 = cfiType_10 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1278 = cfiType_11 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1279 = cfiType_12 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1280 = cfiType_13 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1281 = cfiType_14 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1282 = cfiType_15 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1283 = cfiType_16 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1284 = cfiType_17 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1285 = cfiType_18 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1286 = cfiType_19 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1287 = cfiType_20 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1288 = cfiType_21 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1289 = cfiType_22 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1290 = cfiType_23 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1291 = cfiType_24 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1292 = cfiType_25 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1293 = cfiType_26 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1294 = cfiType_27 == 2'h3; // @[BTB.scala 314:42]
  assign _T_1300 = {_T_1273,_T_1272,_T_1271,_T_1270,_T_1269,_T_1268,_T_1267}; // @[Cat.scala 30:58]
  assign _T_1307 = {_T_1280,_T_1279,_T_1278,_T_1277,_T_1276,_T_1275,_T_1274,_T_1300}; // @[Cat.scala 30:58]
  assign _T_1313 = {_T_1287,_T_1286,_T_1285,_T_1284,_T_1283,_T_1282,_T_1281}; // @[Cat.scala 30:58]
  assign _T_1321 = {_T_1294,_T_1293,_T_1292,_T_1291,_T_1290,_T_1289,_T_1288,_T_1313,_T_1307}; // @[Cat.scala 30:58]
  assign _T_1322 = idxHit & _T_1321; // @[BTB.scala 314:26]
  assign _T_1323 = _T_1322 != 28'h0; // @[BTB.scala 314:67]
  assign _T_1324 = _T_1252 == 3'h0; // @[BTB.scala 55:29]
  assign _GEN_399 = 3'h1 == _T_1254 ? _T_1258_1 : _T_1258_0; // @[BTB.scala 316:22]
  assign _GEN_400 = 3'h2 == _T_1254 ? _T_1258_2 : _GEN_399; // @[BTB.scala 316:22]
  assign _GEN_401 = 3'h3 == _T_1254 ? _T_1258_3 : _GEN_400; // @[BTB.scala 316:22]
  assign _GEN_402 = 3'h4 == _T_1254 ? _T_1258_4 : _GEN_401; // @[BTB.scala 316:22]
  assign _GEN_403 = 3'h5 == _T_1254 ? _T_1258_5 : _GEN_402; // @[BTB.scala 316:22]
  assign _T_1329 = ~_T_1324 & _T_1323; // @[BTB.scala 317:24]
  assign _T_1331 = io_ras_update_bits_cfiType == 2'h2; // @[BTB.scala 321:40]
  assign _T_1332 = _T_1252 < 3'h6; // @[BTB.scala 44:17]
  assign _T_1334 = _T_1252 + 3'h1; // @[BTB.scala 44:42]
  assign _T_1335 = _T_1254 < 3'h5; // @[BTB.scala 45:49]
  assign _T_1338 = _T_1254 + 3'h1; // @[BTB.scala 45:62]
  assign _T_1339 = _T_1335 ? _T_1338 : 3'h0; // @[BTB.scala 45:22]
  assign _T_1341 = io_ras_update_bits_cfiType == 2'h3; // @[BTB.scala 323:46]
  assign _T_1346 = _T_1252 - 3'h1; // @[BTB.scala 51:20]
  assign _T_1347 = _T_1254 > 3'h0; // @[BTB.scala 52:42]
  assign _T_1351 = _T_1254 - 3'h1; // @[BTB.scala 52:50]
  assign io_resp_valid = _T_589[0]; // @[BTB.scala 275:17]
  assign io_resp_bits_taken = _T_1250 ? 1'h0 : 1'h1; // @[BTB.scala 276:22 BTB.scala 308:56]
  assign io_resp_bits_bridx = _T_869 | _T_843; // @[BTB.scala 279:22]
  assign io_resp_bits_target = _T_1329 ? _GEN_403 : _T_765; // @[BTB.scala 277:23 BTB.scala 318:27]
  assign io_resp_bits_entry = {_T_768,_T_785}; // @[BTB.scala 278:22]
  assign io_resp_bits_bht_history = _T_1163; // @[BTB.scala 309:22]
  assign io_resp_bits_bht_value = _T_1161__T_1232_data; // @[BTB.scala 309:22]
  assign io_ras_head_valid = ~_T_1324; // @[BTB.scala 315:23]
  assign io_ras_head_bits = 3'h5 == _T_1254 ? _T_1258_5 : _GEN_402; // @[BTB.scala 316:22]
  assign BTB_cov_read_addr = BTB_state;
  assign BTB_cov_read_data = BTB_cov[BTB_cov_read_addr]; // @[Coverage map for BTB]
  assign BTB_cov_write_data = 1'h1;
  assign BTB_cov_write_addr = BTB_state;
  assign BTB_cov_write_mask = 1'h1;
  assign BTB_cov_write_en = 1'h1;
  assign mux_cond_0 = idxHit[2];
  assign mux_cond_1 = idxHit[16];
  assign mux_cond_2 = idxHit[22];
  assign mux_cond_3 = idxHit[15];
  assign mux_cond_4 = idxHit[0];
  assign mux_cond_5 = idxHit[10];
  assign mux_cond_6 = idxHit[6];
  assign mux_cond_7 = idxHit[5];
  assign mux_cond_8 = idxHit[25];
  assign mux_cond_9 = idxHit[24];
  assign mux_cond_10 = idxHit[11];
  assign mux_cond_11 = idxHit[7];
  assign mux_cond_12 = idxHit[1];
  assign mux_cond_13 = idxHit[27];
  assign mux_cond_14 = idxHit[20];
  assign mux_cond_15 = idxHit[17];
  assign mux_cond_16 = idxHit[18];
  assign mux_cond_17 = idxHit[8];
  assign mux_cond_18 = idxHit[12];
  assign mux_cond_19 = idxHit[3];
  assign mux_cond_20 = idxHit[23];
  assign mux_cond_21 = idxHit[13];
  assign mux_cond_22 = idxHit[21];
  assign mux_cond_23 = idxHit[14];
  assign mux_cond_24 = _T_1156;
  assign mux_cond_25 = idxHit[9];
  assign mux_cond_26 = idxHit[4];
  assign mux_cond_27 = idxHit[19];
  assign mux_cond_28 = idxHit[26];
  assign r_resp_bits_taken_shl = {r_resp_bits_taken, 5'h0};
  assign r_resp_bits_taken_pad = {14'h0,r_resp_bits_taken_shl};
  assign _T_1252_shl = {_T_1252, 7'h0};
  assign _T_1252_pad = {10'h0,_T_1252_shl};
  assign pageValid_shl = {pageValid, 3'h0};
  assign pageValid_pad = {11'h0,pageValid_shl};
  assign r_btb_update_valid_shl = {r_btb_update_valid, 5'h0};
  assign r_btb_update_valid_pad = {14'h0,r_btb_update_valid_shl};
  assign _T_1254_shl = {_T_1254, 3'h0};
  assign _T_1254_pad = {14'h0,_T_1254_shl};
  assign r_resp_valid_shl = {r_resp_valid, 6'h0};
  assign r_resp_valid_pad = {13'h0,r_resp_valid_shl};
  assign r_btb_update_bits_isValid_shl = {r_btb_update_bits_isValid, 11'h0};
  assign r_btb_update_bits_isValid_pad = {8'h0,r_btb_update_bits_isValid_shl};
  assign nextPageRepl_shl = {nextPageRepl, 5'h0};
  assign nextPageRepl_pad = {12'h0,nextPageRepl_shl};
  assign mux_cond_0_shl = {mux_cond_0, 18'h0};
  assign mux_cond_0_pad = {1'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 8'h0};
  assign mux_cond_1_pad = {11'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 15'h0};
  assign mux_cond_2_pad = {4'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 8'h0};
  assign mux_cond_3_pad = {11'h0,mux_cond_3_shl};
  assign mux_cond_4_shl = {mux_cond_4, 1'h0};
  assign mux_cond_4_pad = {18'h0,mux_cond_4_shl};
  assign mux_cond_5_shl = {mux_cond_5, 11'h0};
  assign mux_cond_5_pad = {8'h0,mux_cond_5_shl};
  assign mux_cond_6_shl = {mux_cond_6, 4'h0};
  assign mux_cond_6_pad = {15'h0,mux_cond_6_shl};
  assign mux_cond_7_shl = {mux_cond_7, 15'h0};
  assign mux_cond_7_pad = {4'h0,mux_cond_7_shl};
  assign mux_cond_8_shl = {mux_cond_8, 19'h0};
  assign mux_cond_8_pad = mux_cond_8_shl;
  assign mux_cond_9_shl = {mux_cond_9, 10'h0};
  assign mux_cond_9_pad = {9'h0,mux_cond_9_shl};
  assign mux_cond_10_shl = {mux_cond_10, 6'h0};
  assign mux_cond_10_pad = {13'h0,mux_cond_10_shl};
  assign mux_cond_11_shl = {mux_cond_11, 4'h0};
  assign mux_cond_11_pad = {15'h0,mux_cond_11_shl};
  assign mux_cond_12_shl = {mux_cond_12, 14'h0};
  assign mux_cond_12_pad = {5'h0,mux_cond_12_shl};
  assign mux_cond_13_shl = {mux_cond_13, 3'h0};
  assign mux_cond_13_pad = {16'h0,mux_cond_13_shl};
  assign mux_cond_14_shl = {mux_cond_14, 17'h0};
  assign mux_cond_14_pad = {2'h0,mux_cond_14_shl};
  assign mux_cond_15_shl = {mux_cond_15, 10'h0};
  assign mux_cond_15_pad = {9'h0,mux_cond_15_shl};
  assign mux_cond_16_shl = {mux_cond_16, 18'h0};
  assign mux_cond_16_pad = {1'h0,mux_cond_16_shl};
  assign mux_cond_17_shl = {mux_cond_17, 17'h0};
  assign mux_cond_17_pad = {2'h0,mux_cond_17_shl};
  assign mux_cond_18_shl = {mux_cond_18, 8'h0};
  assign mux_cond_18_pad = {11'h0,mux_cond_18_shl};
  assign mux_cond_19_shl = {mux_cond_19, 8'h0};
  assign mux_cond_19_pad = {11'h0,mux_cond_19_shl};
  assign mux_cond_20_shl = {mux_cond_20, 3'h0};
  assign mux_cond_20_pad = {16'h0,mux_cond_20_shl};
  assign mux_cond_21_shl = {mux_cond_21, 6'h0};
  assign mux_cond_21_pad = {13'h0,mux_cond_21_shl};
  assign mux_cond_22_shl = {mux_cond_22, 19'h0};
  assign mux_cond_22_pad = mux_cond_22_shl;
  assign mux_cond_23_shl = {mux_cond_23, 10'h0};
  assign mux_cond_23_pad = {9'h0,mux_cond_23_shl};
  assign mux_cond_24_shl = {mux_cond_24, 1'h0};
  assign mux_cond_24_pad = {18'h0,mux_cond_24_shl};
  assign mux_cond_25_shl = mux_cond_25;
  assign mux_cond_25_pad = {19'h0,mux_cond_25_shl};
  assign mux_cond_26_shl = {mux_cond_26, 8'h0};
  assign mux_cond_26_pad = {11'h0,mux_cond_26_shl};
  assign mux_cond_27_shl = {mux_cond_27, 2'h0};
  assign mux_cond_27_pad = {17'h0,mux_cond_27_shl};
  assign mux_cond_28_shl = {mux_cond_28, 3'h0};
  assign mux_cond_28_pad = {16'h0,mux_cond_28_shl};
  assign cfiType_4_shl = {cfiType_4, 10'h0};
  assign cfiType_4_pad = {8'h0,cfiType_4_shl};
  assign tgtPages_20_shl = {tgtPages_20, 5'h0};
  assign tgtPages_20_pad = {12'h0,tgtPages_20_shl};
  assign tgtPages_17_shl = {tgtPages_17, 5'h0};
  assign tgtPages_17_pad = {12'h0,tgtPages_17_shl};
  assign tgtPages_3_shl = {tgtPages_3, 5'h0};
  assign tgtPages_3_pad = {12'h0,tgtPages_3_shl};
  assign cfiType_1_shl = {cfiType_1, 10'h0};
  assign cfiType_1_pad = {8'h0,cfiType_1_shl};
  assign tgtPages_2_shl = {tgtPages_2, 5'h0};
  assign tgtPages_2_pad = {12'h0,tgtPages_2_shl};
  assign cfiType_18_shl = {cfiType_18, 10'h0};
  assign cfiType_18_pad = {8'h0,cfiType_18_shl};
  assign tgtPages_26_shl = {tgtPages_26, 5'h0};
  assign tgtPages_26_pad = {12'h0,tgtPages_26_shl};
  assign cfiType_20_shl = {cfiType_20, 10'h0};
  assign cfiType_20_pad = {8'h0,cfiType_20_shl};
  assign cfiType_22_shl = {cfiType_22, 10'h0};
  assign cfiType_22_pad = {8'h0,cfiType_22_shl};
  assign cfiType_23_shl = {cfiType_23, 10'h0};
  assign cfiType_23_pad = {8'h0,cfiType_23_shl};
  assign cfiType_0_shl = {cfiType_0, 10'h0};
  assign cfiType_0_pad = {8'h0,cfiType_0_shl};
  assign tgtPages_11_shl = {tgtPages_11, 5'h0};
  assign tgtPages_11_pad = {12'h0,tgtPages_11_shl};
  assign cfiType_7_shl = {cfiType_7, 10'h0};
  assign cfiType_7_pad = {8'h0,cfiType_7_shl};
  assign cfiType_19_shl = {cfiType_19, 10'h0};
  assign cfiType_19_pad = {8'h0,cfiType_19_shl};
  assign cfiType_17_shl = {cfiType_17, 10'h0};
  assign cfiType_17_pad = {8'h0,cfiType_17_shl};
  assign cfiType_25_shl = {cfiType_25, 10'h0};
  assign cfiType_25_pad = {8'h0,cfiType_25_shl};
  assign cfiType_3_shl = {cfiType_3, 10'h0};
  assign cfiType_3_pad = {8'h0,cfiType_3_shl};
  assign cfiType_10_shl = {cfiType_10, 10'h0};
  assign cfiType_10_pad = {8'h0,cfiType_10_shl};
  assign tgtPages_14_shl = {tgtPages_14, 5'h0};
  assign tgtPages_14_pad = {12'h0,tgtPages_14_shl};
  assign cfiType_2_shl = {cfiType_2, 10'h0};
  assign cfiType_2_pad = {8'h0,cfiType_2_shl};
  assign cfiType_16_shl = {cfiType_16, 10'h0};
  assign cfiType_16_pad = {8'h0,cfiType_16_shl};
  assign tgtPages_0_shl = {tgtPages_0, 5'h0};
  assign tgtPages_0_pad = {12'h0,tgtPages_0_shl};
  assign tgtPages_21_shl = {tgtPages_21, 5'h0};
  assign tgtPages_21_pad = {12'h0,tgtPages_21_shl};
  assign tgtPages_5_shl = {tgtPages_5, 5'h0};
  assign tgtPages_5_pad = {12'h0,tgtPages_5_shl};
  assign tgtPages_4_shl = {tgtPages_4, 5'h0};
  assign tgtPages_4_pad = {12'h0,tgtPages_4_shl};
  assign cfiType_9_shl = {cfiType_9, 10'h0};
  assign cfiType_9_pad = {8'h0,cfiType_9_shl};
  assign tgtPages_25_shl = {tgtPages_25, 5'h0};
  assign tgtPages_25_pad = {12'h0,tgtPages_25_shl};
  assign cfiType_8_shl = {cfiType_8, 10'h0};
  assign cfiType_8_pad = {8'h0,cfiType_8_shl};
  assign tgtPages_24_shl = {tgtPages_24, 5'h0};
  assign tgtPages_24_pad = {12'h0,tgtPages_24_shl};
  assign cfiType_26_shl = {cfiType_26, 10'h0};
  assign cfiType_26_pad = {8'h0,cfiType_26_shl};
  assign tgtPages_13_shl = {tgtPages_13, 5'h0};
  assign tgtPages_13_pad = {12'h0,tgtPages_13_shl};
  assign cfiType_14_shl = {cfiType_14, 10'h0};
  assign cfiType_14_pad = {8'h0,cfiType_14_shl};
  assign cfiType_11_shl = {cfiType_11, 10'h0};
  assign cfiType_11_pad = {8'h0,cfiType_11_shl};
  assign tgtPages_16_shl = {tgtPages_16, 5'h0};
  assign tgtPages_16_pad = {12'h0,tgtPages_16_shl};
  assign cfiType_15_shl = {cfiType_15, 10'h0};
  assign cfiType_15_pad = {8'h0,cfiType_15_shl};
  assign cfiType_24_shl = {cfiType_24, 10'h0};
  assign cfiType_24_pad = {8'h0,cfiType_24_shl};
  assign tgtPages_18_shl = {tgtPages_18, 5'h0};
  assign tgtPages_18_pad = {12'h0,tgtPages_18_shl};
  assign cfiType_21_shl = {cfiType_21, 10'h0};
  assign cfiType_21_pad = {8'h0,cfiType_21_shl};
  assign tgtPages_12_shl = {tgtPages_12, 5'h0};
  assign tgtPages_12_pad = {12'h0,tgtPages_12_shl};
  assign tgtPages_10_shl = {tgtPages_10, 5'h0};
  assign tgtPages_10_pad = {12'h0,tgtPages_10_shl};
  assign tgtPages_15_shl = {tgtPages_15, 5'h0};
  assign tgtPages_15_pad = {12'h0,tgtPages_15_shl};
  assign tgtPages_22_shl = {tgtPages_22, 5'h0};
  assign tgtPages_22_pad = {12'h0,tgtPages_22_shl};
  assign tgtPages_19_shl = {tgtPages_19, 5'h0};
  assign tgtPages_19_pad = {12'h0,tgtPages_19_shl};
  assign cfiType_13_shl = {cfiType_13, 10'h0};
  assign cfiType_13_pad = {8'h0,cfiType_13_shl};
  assign cfiType_6_shl = {cfiType_6, 10'h0};
  assign cfiType_6_pad = {8'h0,cfiType_6_shl};
  assign tgtPages_6_shl = {tgtPages_6, 5'h0};
  assign tgtPages_6_pad = {12'h0,tgtPages_6_shl};
  assign cfiType_27_shl = {cfiType_27, 10'h0};
  assign cfiType_27_pad = {8'h0,cfiType_27_shl};
  assign tgtPages_23_shl = {tgtPages_23, 5'h0};
  assign tgtPages_23_pad = {12'h0,tgtPages_23_shl};
  assign cfiType_12_shl = {cfiType_12, 10'h0};
  assign cfiType_12_pad = {8'h0,cfiType_12_shl};
  assign tgtPages_8_shl = {tgtPages_8, 5'h0};
  assign tgtPages_8_pad = {12'h0,tgtPages_8_shl};
  assign tgtPages_1_shl = {tgtPages_1, 5'h0};
  assign tgtPages_1_pad = {12'h0,tgtPages_1_shl};
  assign tgtPages_9_shl = {tgtPages_9, 5'h0};
  assign tgtPages_9_pad = {12'h0,tgtPages_9_shl};
  assign cfiType_5_shl = {cfiType_5, 10'h0};
  assign cfiType_5_pad = {8'h0,cfiType_5_shl};
  assign tgtPages_7_shl = {tgtPages_7, 5'h0};
  assign tgtPages_7_pad = {12'h0,tgtPages_7_shl};
  assign tgtPages_27_shl = {tgtPages_27, 5'h0};
  assign tgtPages_27_pad = {12'h0,tgtPages_27_shl};
  assign BTB_xor31 = r_resp_bits_taken_pad ^ _T_1252_pad;
  assign BTB_xor66 = r_btb_update_valid_pad ^ _T_1254_pad;
  assign BTB_xor32 = pageValid_pad ^ BTB_xor66;
  assign BTB_xor15 = BTB_xor31 ^ BTB_xor32;
  assign BTB_xor68 = r_btb_update_bits_isValid_pad ^ nextPageRepl_pad;
  assign BTB_xor33 = r_resp_valid_pad ^ BTB_xor68;
  assign BTB_xor70 = mux_cond_1_pad ^ mux_cond_2_pad;
  assign BTB_xor34 = mux_cond_0_pad ^ BTB_xor70;
  assign BTB_xor16 = BTB_xor33 ^ BTB_xor34;
  assign BTB_xor7 = BTB_xor15 ^ BTB_xor16;
  assign BTB_xor72 = mux_cond_4_pad ^ mux_cond_5_pad;
  assign BTB_xor35 = mux_cond_3_pad ^ BTB_xor72;
  assign BTB_xor74 = mux_cond_7_pad ^ mux_cond_8_pad;
  assign BTB_xor36 = mux_cond_6_pad ^ BTB_xor74;
  assign BTB_xor17 = BTB_xor35 ^ BTB_xor36;
  assign BTB_xor76 = mux_cond_10_pad ^ mux_cond_11_pad;
  assign BTB_xor37 = mux_cond_9_pad ^ BTB_xor76;
  assign BTB_xor78 = mux_cond_13_pad ^ mux_cond_14_pad;
  assign BTB_xor38 = mux_cond_12_pad ^ BTB_xor78;
  assign BTB_xor18 = BTB_xor37 ^ BTB_xor38;
  assign BTB_xor8 = BTB_xor17 ^ BTB_xor18;
  assign BTB_xor3 = BTB_xor7 ^ BTB_xor8;
  assign BTB_xor39 = mux_cond_15_pad ^ mux_cond_16_pad;
  assign BTB_xor82 = mux_cond_18_pad ^ mux_cond_19_pad;
  assign BTB_xor40 = mux_cond_17_pad ^ BTB_xor82;
  assign BTB_xor19 = BTB_xor39 ^ BTB_xor40;
  assign BTB_xor84 = mux_cond_21_pad ^ mux_cond_22_pad;
  assign BTB_xor41 = mux_cond_20_pad ^ BTB_xor84;
  assign BTB_xor86 = mux_cond_24_pad ^ mux_cond_25_pad;
  assign BTB_xor42 = mux_cond_23_pad ^ BTB_xor86;
  assign BTB_xor20 = BTB_xor41 ^ BTB_xor42;
  assign BTB_xor9 = BTB_xor19 ^ BTB_xor20;
  assign BTB_xor88 = mux_cond_27_pad ^ mux_cond_28_pad;
  assign BTB_xor43 = mux_cond_26_pad ^ BTB_xor88;
  assign BTB_xor90 = tgtPages_20_pad ^ tgtPages_17_pad;
  assign BTB_xor44 = cfiType_4_pad ^ BTB_xor90;
  assign BTB_xor21 = BTB_xor43 ^ BTB_xor44;
  assign BTB_xor92 = cfiType_1_pad ^ tgtPages_2_pad;
  assign BTB_xor45 = tgtPages_3_pad ^ BTB_xor92;
  assign BTB_xor94 = tgtPages_26_pad ^ cfiType_20_pad;
  assign BTB_xor46 = cfiType_18_pad ^ BTB_xor94;
  assign BTB_xor22 = BTB_xor45 ^ BTB_xor46;
  assign BTB_xor10 = BTB_xor21 ^ BTB_xor22;
  assign BTB_xor4 = BTB_xor9 ^ BTB_xor10;
  assign BTB_xor1 = BTB_xor3 ^ BTB_xor4;
  assign BTB_xor47 = cfiType_22_pad ^ cfiType_23_pad;
  assign BTB_xor98 = tgtPages_11_pad ^ cfiType_7_pad;
  assign BTB_xor48 = cfiType_0_pad ^ BTB_xor98;
  assign BTB_xor23 = BTB_xor47 ^ BTB_xor48;
  assign BTB_xor100 = cfiType_17_pad ^ cfiType_25_pad;
  assign BTB_xor49 = cfiType_19_pad ^ BTB_xor100;
  assign BTB_xor102 = cfiType_10_pad ^ tgtPages_14_pad;
  assign BTB_xor50 = cfiType_3_pad ^ BTB_xor102;
  assign BTB_xor24 = BTB_xor49 ^ BTB_xor50;
  assign BTB_xor11 = BTB_xor23 ^ BTB_xor24;
  assign BTB_xor104 = cfiType_16_pad ^ tgtPages_0_pad;
  assign BTB_xor51 = cfiType_2_pad ^ BTB_xor104;
  assign BTB_xor106 = tgtPages_5_pad ^ tgtPages_4_pad;
  assign BTB_xor52 = tgtPages_21_pad ^ BTB_xor106;
  assign BTB_xor25 = BTB_xor51 ^ BTB_xor52;
  assign BTB_xor108 = tgtPages_25_pad ^ cfiType_8_pad;
  assign BTB_xor53 = cfiType_9_pad ^ BTB_xor108;
  assign BTB_xor110 = cfiType_26_pad ^ tgtPages_13_pad;
  assign BTB_xor54 = tgtPages_24_pad ^ BTB_xor110;
  assign BTB_xor26 = BTB_xor53 ^ BTB_xor54;
  assign BTB_xor12 = BTB_xor25 ^ BTB_xor26;
  assign BTB_xor5 = BTB_xor11 ^ BTB_xor12;
  assign BTB_xor112 = cfiType_11_pad ^ tgtPages_16_pad;
  assign BTB_xor55 = cfiType_14_pad ^ BTB_xor112;
  assign BTB_xor114 = cfiType_24_pad ^ tgtPages_18_pad;
  assign BTB_xor56 = cfiType_15_pad ^ BTB_xor114;
  assign BTB_xor27 = BTB_xor55 ^ BTB_xor56;
  assign BTB_xor116 = tgtPages_12_pad ^ tgtPages_10_pad;
  assign BTB_xor57 = cfiType_21_pad ^ BTB_xor116;
  assign BTB_xor118 = tgtPages_22_pad ^ tgtPages_19_pad;
  assign BTB_xor58 = tgtPages_15_pad ^ BTB_xor118;
  assign BTB_xor28 = BTB_xor57 ^ BTB_xor58;
  assign BTB_xor13 = BTB_xor27 ^ BTB_xor28;
  assign BTB_xor120 = cfiType_6_pad ^ tgtPages_6_pad;
  assign BTB_xor59 = cfiType_13_pad ^ BTB_xor120;
  assign BTB_xor122 = tgtPages_23_pad ^ cfiType_12_pad;
  assign BTB_xor60 = cfiType_27_pad ^ BTB_xor122;
  assign BTB_xor29 = BTB_xor59 ^ BTB_xor60;
  assign BTB_xor124 = tgtPages_1_pad ^ tgtPages_9_pad;
  assign BTB_xor61 = tgtPages_8_pad ^ BTB_xor124;
  assign BTB_xor126 = tgtPages_7_pad ^ tgtPages_27_pad;
  assign BTB_xor62 = cfiType_5_pad ^ BTB_xor126;
  assign BTB_xor30 = BTB_xor61 ^ BTB_xor62;
  assign BTB_xor14 = BTB_xor29 ^ BTB_xor30;
  assign BTB_xor6 = BTB_xor13 ^ BTB_xor14;
  assign BTB_xor2 = BTB_xor5 ^ BTB_xor6;
  assign BTB_xor0 = BTB_xor1 ^ BTB_xor2;
  assign io_covSum = BTB_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    _T_1161[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  idxs_0 = _RAND_1[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  idxs_1 = _RAND_2[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  idxs_2 = _RAND_3[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  idxs_3 = _RAND_4[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  idxs_4 = _RAND_5[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  idxs_5 = _RAND_6[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  idxs_6 = _RAND_7[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  idxs_7 = _RAND_8[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idxs_8 = _RAND_9[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idxs_9 = _RAND_10[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  idxs_10 = _RAND_11[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  idxs_11 = _RAND_12[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  idxs_12 = _RAND_13[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  idxs_13 = _RAND_14[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  idxs_14 = _RAND_15[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  idxs_15 = _RAND_16[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  idxs_16 = _RAND_17[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  idxs_17 = _RAND_18[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  idxs_18 = _RAND_19[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  idxs_19 = _RAND_20[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  idxs_20 = _RAND_21[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  idxs_21 = _RAND_22[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  idxs_22 = _RAND_23[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  idxs_23 = _RAND_24[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  idxs_24 = _RAND_25[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  idxs_25 = _RAND_26[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  idxs_26 = _RAND_27[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  idxs_27 = _RAND_28[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  idxPages_0 = _RAND_29[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  idxPages_1 = _RAND_30[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  idxPages_2 = _RAND_31[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  idxPages_3 = _RAND_32[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  idxPages_4 = _RAND_33[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  idxPages_5 = _RAND_34[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  idxPages_6 = _RAND_35[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  idxPages_7 = _RAND_36[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  idxPages_8 = _RAND_37[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  idxPages_9 = _RAND_38[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  idxPages_10 = _RAND_39[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  idxPages_11 = _RAND_40[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  idxPages_12 = _RAND_41[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  idxPages_13 = _RAND_42[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  idxPages_14 = _RAND_43[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  idxPages_15 = _RAND_44[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  idxPages_16 = _RAND_45[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  idxPages_17 = _RAND_46[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  idxPages_18 = _RAND_47[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  idxPages_19 = _RAND_48[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  idxPages_20 = _RAND_49[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  idxPages_21 = _RAND_50[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  idxPages_22 = _RAND_51[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  idxPages_23 = _RAND_52[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  idxPages_24 = _RAND_53[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  idxPages_25 = _RAND_54[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  idxPages_26 = _RAND_55[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  idxPages_27 = _RAND_56[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  tgts_0 = _RAND_57[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  tgts_1 = _RAND_58[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  tgts_2 = _RAND_59[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  tgts_3 = _RAND_60[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  tgts_4 = _RAND_61[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  tgts_5 = _RAND_62[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  tgts_6 = _RAND_63[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  tgts_7 = _RAND_64[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  tgts_8 = _RAND_65[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  tgts_9 = _RAND_66[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  tgts_10 = _RAND_67[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  tgts_11 = _RAND_68[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  tgts_12 = _RAND_69[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  tgts_13 = _RAND_70[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  tgts_14 = _RAND_71[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  tgts_15 = _RAND_72[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  tgts_16 = _RAND_73[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  tgts_17 = _RAND_74[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  tgts_18 = _RAND_75[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  tgts_19 = _RAND_76[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  tgts_20 = _RAND_77[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  tgts_21 = _RAND_78[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  tgts_22 = _RAND_79[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  tgts_23 = _RAND_80[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  tgts_24 = _RAND_81[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  tgts_25 = _RAND_82[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  tgts_26 = _RAND_83[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  tgts_27 = _RAND_84[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  tgtPages_0 = _RAND_85[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  tgtPages_1 = _RAND_86[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  tgtPages_2 = _RAND_87[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  tgtPages_3 = _RAND_88[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  tgtPages_4 = _RAND_89[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  tgtPages_5 = _RAND_90[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  tgtPages_6 = _RAND_91[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  tgtPages_7 = _RAND_92[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  tgtPages_8 = _RAND_93[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  tgtPages_9 = _RAND_94[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  tgtPages_10 = _RAND_95[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  tgtPages_11 = _RAND_96[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  tgtPages_12 = _RAND_97[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  tgtPages_13 = _RAND_98[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  tgtPages_14 = _RAND_99[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  tgtPages_15 = _RAND_100[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  tgtPages_16 = _RAND_101[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  tgtPages_17 = _RAND_102[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  tgtPages_18 = _RAND_103[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  tgtPages_19 = _RAND_104[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  tgtPages_20 = _RAND_105[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  tgtPages_21 = _RAND_106[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  tgtPages_22 = _RAND_107[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  tgtPages_23 = _RAND_108[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  tgtPages_24 = _RAND_109[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  tgtPages_25 = _RAND_110[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  tgtPages_26 = _RAND_111[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  tgtPages_27 = _RAND_112[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  pages_0 = _RAND_113[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  pages_1 = _RAND_114[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  pages_2 = _RAND_115[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  pages_3 = _RAND_116[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  pages_4 = _RAND_117[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  pages_5 = _RAND_118[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  pageValid = _RAND_119[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  isValid = _RAND_120[27:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  cfiType_0 = _RAND_121[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  cfiType_1 = _RAND_122[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  cfiType_2 = _RAND_123[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  cfiType_3 = _RAND_124[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  cfiType_4 = _RAND_125[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  cfiType_5 = _RAND_126[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  cfiType_6 = _RAND_127[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  cfiType_7 = _RAND_128[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  cfiType_8 = _RAND_129[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  cfiType_9 = _RAND_130[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  cfiType_10 = _RAND_131[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  cfiType_11 = _RAND_132[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  cfiType_12 = _RAND_133[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  cfiType_13 = _RAND_134[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  cfiType_14 = _RAND_135[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  cfiType_15 = _RAND_136[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  cfiType_16 = _RAND_137[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  cfiType_17 = _RAND_138[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  cfiType_18 = _RAND_139[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  cfiType_19 = _RAND_140[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  cfiType_20 = _RAND_141[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  cfiType_21 = _RAND_142[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  cfiType_22 = _RAND_143[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  cfiType_23 = _RAND_144[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  cfiType_24 = _RAND_145[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  cfiType_25 = _RAND_146[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  cfiType_26 = _RAND_147[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  cfiType_27 = _RAND_148[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  brIdx_0 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  brIdx_1 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  brIdx_2 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  brIdx_3 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  brIdx_4 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  brIdx_5 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  brIdx_6 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  brIdx_7 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  brIdx_8 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  brIdx_9 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  brIdx_10 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  brIdx_11 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  brIdx_12 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  brIdx_13 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  brIdx_14 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  brIdx_15 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  brIdx_16 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  brIdx_17 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  brIdx_18 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  brIdx_19 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  brIdx_20 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  brIdx_21 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  brIdx_22 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  brIdx_23 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  brIdx_24 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  brIdx_25 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  brIdx_26 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  brIdx_27 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  r_btb_update_valid = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  r_btb_update_bits_prediction_entry = _RAND_178[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {2{`RANDOM}};
  r_btb_update_bits_pc = _RAND_179[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  r_btb_update_bits_isValid = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {2{`RANDOM}};
  r_btb_update_bits_br_pc = _RAND_181[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  r_btb_update_bits_cfiType = _RAND_182[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  nextPageRepl = _RAND_183[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_373 = _RAND_184[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  r_resp_valid = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  r_resp_bits_taken = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  r_resp_bits_entry = _RAND_187[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_1163 = _RAND_188[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_1252 = _RAND_189[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_1254 = _RAND_190[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {2{`RANDOM}};
  _T_1258_0 = _RAND_191[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {2{`RANDOM}};
  _T_1258_1 = _RAND_192[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {2{`RANDOM}};
  _T_1258_2 = _RAND_193[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {2{`RANDOM}};
  _T_1258_3 = _RAND_194[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {2{`RANDOM}};
  _T_1258_4 = _RAND_195[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {2{`RANDOM}};
  _T_1258_5 = _RAND_196[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  BTB_state = _RAND_197[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    BTB_cov[initvar] = _RAND_198[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  BTB_covSum = _RAND_199[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_1161__T_1245_en & _T_1161__T_1245_mask) begin
      _T_1161[_T_1161__T_1245_addr] <= _T_1161__T_1245_data; // @[BTB.scala 113:26]
    end
    if (metaReset) begin
      idxs_0 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h0 == waddr) begin
        idxs_0 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_1 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h1 == waddr) begin
        idxs_1 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_2 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h2 == waddr) begin
        idxs_2 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_3 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h3 == waddr) begin
        idxs_3 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_4 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h4 == waddr) begin
        idxs_4 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_5 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h5 == waddr) begin
        idxs_5 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_6 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h6 == waddr) begin
        idxs_6 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_7 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h7 == waddr) begin
        idxs_7 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_8 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h8 == waddr) begin
        idxs_8 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_9 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h9 == waddr) begin
        idxs_9 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_10 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'ha == waddr) begin
        idxs_10 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_11 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'hb == waddr) begin
        idxs_11 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_12 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'hc == waddr) begin
        idxs_12 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_13 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'hd == waddr) begin
        idxs_13 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_14 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'he == waddr) begin
        idxs_14 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_15 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'hf == waddr) begin
        idxs_15 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_16 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h10 == waddr) begin
        idxs_16 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_17 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h11 == waddr) begin
        idxs_17 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_18 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h12 == waddr) begin
        idxs_18 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_19 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h13 == waddr) begin
        idxs_19 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_20 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h14 == waddr) begin
        idxs_20 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_21 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h15 == waddr) begin
        idxs_21 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_22 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h16 == waddr) begin
        idxs_22 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_23 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h17 == waddr) begin
        idxs_23 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_24 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h18 == waddr) begin
        idxs_24 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_25 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h19 == waddr) begin
        idxs_25 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_26 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h1a == waddr) begin
        idxs_26 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_27 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h1b == waddr) begin
        idxs_27 <= r_btb_update_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxPages_0 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h0 == waddr) begin
        idxPages_0 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_1 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h1 == waddr) begin
        idxPages_1 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_2 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h2 == waddr) begin
        idxPages_2 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_3 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h3 == waddr) begin
        idxPages_3 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_4 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h4 == waddr) begin
        idxPages_4 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_5 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h5 == waddr) begin
        idxPages_5 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_6 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h6 == waddr) begin
        idxPages_6 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_7 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h7 == waddr) begin
        idxPages_7 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_8 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h8 == waddr) begin
        idxPages_8 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_9 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h9 == waddr) begin
        idxPages_9 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_10 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'ha == waddr) begin
        idxPages_10 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_11 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'hb == waddr) begin
        idxPages_11 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_12 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'hc == waddr) begin
        idxPages_12 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_13 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'hd == waddr) begin
        idxPages_13 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_14 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'he == waddr) begin
        idxPages_14 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_15 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'hf == waddr) begin
        idxPages_15 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_16 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h10 == waddr) begin
        idxPages_16 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_17 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h11 == waddr) begin
        idxPages_17 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_18 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h12 == waddr) begin
        idxPages_18 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_19 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h13 == waddr) begin
        idxPages_19 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_20 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h14 == waddr) begin
        idxPages_20 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_21 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h15 == waddr) begin
        idxPages_21 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_22 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h16 == waddr) begin
        idxPages_22 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_23 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h17 == waddr) begin
        idxPages_23 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_24 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h18 == waddr) begin
        idxPages_24 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_25 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h19 == waddr) begin
        idxPages_25 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_26 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h1a == waddr) begin
        idxPages_26 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      idxPages_27 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h1b == waddr) begin
        idxPages_27 <= _T_475[2:0];
      end
    end
    if (metaReset) begin
      tgts_0 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h0 == waddr) begin
        tgts_0 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_1 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h1 == waddr) begin
        tgts_1 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_2 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h2 == waddr) begin
        tgts_2 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_3 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h3 == waddr) begin
        tgts_3 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_4 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h4 == waddr) begin
        tgts_4 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_5 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h5 == waddr) begin
        tgts_5 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_6 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h6 == waddr) begin
        tgts_6 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_7 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h7 == waddr) begin
        tgts_7 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_8 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h8 == waddr) begin
        tgts_8 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_9 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h9 == waddr) begin
        tgts_9 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_10 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'ha == waddr) begin
        tgts_10 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_11 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'hb == waddr) begin
        tgts_11 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_12 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'hc == waddr) begin
        tgts_12 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_13 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'hd == waddr) begin
        tgts_13 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_14 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'he == waddr) begin
        tgts_14 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_15 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'hf == waddr) begin
        tgts_15 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_16 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h10 == waddr) begin
        tgts_16 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_17 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h11 == waddr) begin
        tgts_17 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_18 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h12 == waddr) begin
        tgts_18 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_19 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h13 == waddr) begin
        tgts_19 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_20 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h14 == waddr) begin
        tgts_20 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_21 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h15 == waddr) begin
        tgts_21 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_22 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h16 == waddr) begin
        tgts_22 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_23 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h17 == waddr) begin
        tgts_23 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_24 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h18 == waddr) begin
        tgts_24 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_25 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h19 == waddr) begin
        tgts_25 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_26 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h1a == waddr) begin
        tgts_26 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgts_27 <= 13'h0;
    end else if (r_btb_update_valid) begin
      if (5'h1b == waddr) begin
        tgts_27 <= io_req_bits_addr[13:1];
      end
    end
    if (metaReset) begin
      tgtPages_0 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h0 == waddr) begin
        tgtPages_0 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_1 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h1 == waddr) begin
        tgtPages_1 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_2 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h2 == waddr) begin
        tgtPages_2 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_3 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h3 == waddr) begin
        tgtPages_3 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_4 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h4 == waddr) begin
        tgtPages_4 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_5 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h5 == waddr) begin
        tgtPages_5 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_6 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h6 == waddr) begin
        tgtPages_6 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_7 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h7 == waddr) begin
        tgtPages_7 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_8 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h8 == waddr) begin
        tgtPages_8 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_9 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h9 == waddr) begin
        tgtPages_9 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_10 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'ha == waddr) begin
        tgtPages_10 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_11 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'hb == waddr) begin
        tgtPages_11 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_12 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'hc == waddr) begin
        tgtPages_12 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_13 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'hd == waddr) begin
        tgtPages_13 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_14 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'he == waddr) begin
        tgtPages_14 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_15 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'hf == waddr) begin
        tgtPages_15 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_16 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h10 == waddr) begin
        tgtPages_16 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_17 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h11 == waddr) begin
        tgtPages_17 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_18 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h12 == waddr) begin
        tgtPages_18 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_19 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h13 == waddr) begin
        tgtPages_19 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_20 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h14 == waddr) begin
        tgtPages_20 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_21 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h15 == waddr) begin
        tgtPages_21 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_22 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h16 == waddr) begin
        tgtPages_22 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_23 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h17 == waddr) begin
        tgtPages_23 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_24 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h18 == waddr) begin
        tgtPages_24 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_25 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h19 == waddr) begin
        tgtPages_25 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_26 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h1a == waddr) begin
        tgtPages_26 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_27 <= 3'h0;
    end else if (r_btb_update_valid) begin
      if (5'h1b == waddr) begin
        tgtPages_27 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      pages_0 <= 25'h0;
    end else if (r_btb_update_valid) begin
      if (_T_486[0]) begin
        if (~idxPageUpdate[0]) begin
          pages_0 <= r_btb_update_bits_pc[38:14];
        end else begin
          pages_0 <= io_req_bits_addr[38:14];
        end
      end
    end
    if (metaReset) begin
      pages_1 <= 25'h0;
    end else if (r_btb_update_valid) begin
      if (_T_493[1]) begin
        if (~idxPageUpdate[0]) begin
          pages_1 <= io_req_bits_addr[38:14];
        end else begin
          pages_1 <= r_btb_update_bits_pc[38:14];
        end
      end
    end
    if (metaReset) begin
      pages_2 <= 25'h0;
    end else if (r_btb_update_valid) begin
      if (_T_486[2]) begin
        if (~idxPageUpdate[0]) begin
          pages_2 <= r_btb_update_bits_pc[38:14];
        end else begin
          pages_2 <= io_req_bits_addr[38:14];
        end
      end
    end
    if (metaReset) begin
      pages_3 <= 25'h0;
    end else if (r_btb_update_valid) begin
      if (_T_493[3]) begin
        if (~idxPageUpdate[0]) begin
          pages_3 <= io_req_bits_addr[38:14];
        end else begin
          pages_3 <= r_btb_update_bits_pc[38:14];
        end
      end
    end
    if (metaReset) begin
      pages_4 <= 25'h0;
    end else if (r_btb_update_valid) begin
      if (_T_486[4]) begin
        if (~idxPageUpdate[0]) begin
          pages_4 <= r_btb_update_bits_pc[38:14];
        end else begin
          pages_4 <= io_req_bits_addr[38:14];
        end
      end
    end
    if (metaReset) begin
      pages_5 <= 25'h0;
    end else if (r_btb_update_valid) begin
      if (_T_493[5]) begin
        if (~idxPageUpdate[0]) begin
          pages_5 <= io_req_bits_addr[38:14];
        end else begin
          pages_5 <= r_btb_update_bits_pc[38:14];
        end
      end
    end
    if (metaReset) begin
      pageValid <= 6'h0;
    end else if (reset) begin
      pageValid <= 6'h0;
    end else begin
      pageValid <= _GEN_373[5:0];
    end
    if (metaReset) begin
      isValid <= 28'h0;
    end else if (reset) begin
      isValid <= 28'h0;
    end else begin
      isValid <= _GEN_381[27:0];
    end
    if (metaReset) begin
      cfiType_0 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'h0 == waddr) begin
        cfiType_0 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_1 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'h1 == waddr) begin
        cfiType_1 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_2 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'h2 == waddr) begin
        cfiType_2 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_3 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'h3 == waddr) begin
        cfiType_3 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_4 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'h4 == waddr) begin
        cfiType_4 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_5 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'h5 == waddr) begin
        cfiType_5 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_6 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'h6 == waddr) begin
        cfiType_6 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_7 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'h7 == waddr) begin
        cfiType_7 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_8 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'h8 == waddr) begin
        cfiType_8 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_9 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'h9 == waddr) begin
        cfiType_9 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_10 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'ha == waddr) begin
        cfiType_10 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_11 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'hb == waddr) begin
        cfiType_11 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_12 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'hc == waddr) begin
        cfiType_12 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_13 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'hd == waddr) begin
        cfiType_13 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_14 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'he == waddr) begin
        cfiType_14 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_15 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'hf == waddr) begin
        cfiType_15 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_16 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'h10 == waddr) begin
        cfiType_16 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_17 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'h11 == waddr) begin
        cfiType_17 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_18 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'h12 == waddr) begin
        cfiType_18 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_19 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'h13 == waddr) begin
        cfiType_19 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_20 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'h14 == waddr) begin
        cfiType_20 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_21 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'h15 == waddr) begin
        cfiType_21 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_22 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'h16 == waddr) begin
        cfiType_22 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_23 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'h17 == waddr) begin
        cfiType_23 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_24 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'h18 == waddr) begin
        cfiType_24 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_25 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'h19 == waddr) begin
        cfiType_25 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_26 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'h1a == waddr) begin
        cfiType_26 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_27 <= 2'h0;
    end else if (r_btb_update_valid) begin
      if (5'h1b == waddr) begin
        cfiType_27 <= r_btb_update_bits_cfiType;
      end
    end
    if (metaReset) begin
      brIdx_0 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'h0 == waddr) begin
        brIdx_0 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_1 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'h1 == waddr) begin
        brIdx_1 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_2 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'h2 == waddr) begin
        brIdx_2 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_3 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'h3 == waddr) begin
        brIdx_3 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_4 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'h4 == waddr) begin
        brIdx_4 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_5 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'h5 == waddr) begin
        brIdx_5 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_6 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'h6 == waddr) begin
        brIdx_6 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_7 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'h7 == waddr) begin
        brIdx_7 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_8 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'h8 == waddr) begin
        brIdx_8 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_9 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'h9 == waddr) begin
        brIdx_9 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_10 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'ha == waddr) begin
        brIdx_10 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_11 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'hb == waddr) begin
        brIdx_11 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_12 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'hc == waddr) begin
        brIdx_12 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_13 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'hd == waddr) begin
        brIdx_13 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_14 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'he == waddr) begin
        brIdx_14 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_15 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'hf == waddr) begin
        brIdx_15 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_16 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'h10 == waddr) begin
        brIdx_16 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_17 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'h11 == waddr) begin
        brIdx_17 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_18 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'h12 == waddr) begin
        brIdx_18 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_19 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'h13 == waddr) begin
        brIdx_19 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_20 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'h14 == waddr) begin
        brIdx_20 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_21 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'h15 == waddr) begin
        brIdx_21 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_22 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'h16 == waddr) begin
        brIdx_22 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_23 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'h17 == waddr) begin
        brIdx_23 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_24 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'h18 == waddr) begin
        brIdx_24 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_25 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'h19 == waddr) begin
        brIdx_25 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_26 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'h1a == waddr) begin
        brIdx_26 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_27 <= 1'h0;
    end else if (r_btb_update_valid) begin
      if (5'h1b == waddr) begin
        brIdx_27 <= r_btb_update_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      r_btb_update_valid <= 1'h0;
    end else if (reset) begin
      r_btb_update_valid <= 1'h0;
    end else begin
      r_btb_update_valid <= io_btb_update_valid;
    end
    if (metaReset) begin
      r_btb_update_bits_prediction_entry <= 5'h0;
    end else if (io_btb_update_valid) begin
      r_btb_update_bits_prediction_entry <= io_btb_update_bits_prediction_entry;
    end
    if (metaReset) begin
      r_btb_update_bits_pc <= 39'h0;
    end else if (io_btb_update_valid) begin
      r_btb_update_bits_pc <= io_btb_update_bits_pc;
    end
    if (metaReset) begin
      r_btb_update_bits_isValid <= 1'h0;
    end else if (io_btb_update_valid) begin
      r_btb_update_bits_isValid <= io_btb_update_bits_isValid;
    end
    if (metaReset) begin
      r_btb_update_bits_br_pc <= 39'h0;
    end else if (io_btb_update_valid) begin
      r_btb_update_bits_br_pc <= io_btb_update_bits_br_pc;
    end
    if (metaReset) begin
      r_btb_update_bits_cfiType <= 2'h0;
    end else if (io_btb_update_valid) begin
      r_btb_update_bits_cfiType <= io_btb_update_bits_cfiType;
    end
    if (metaReset) begin
      nextPageRepl <= 3'h0;
    end else if (_T_364) begin
      if (_T_369) begin
        nextPageRepl <= {{2'd0}, _T_368[0]};
      end else begin
        nextPageRepl <= _T_368;
      end
    end
    if (metaReset) begin
      _T_373 <= 27'h0;
    end else if (_T_420) begin
      _T_373 <= _T_466[27:1];
    end
    if (metaReset) begin
      r_resp_valid <= 1'h0;
    end else if (reset) begin
      r_resp_valid <= 1'h0;
    end else begin
      r_resp_valid <= io_resp_valid;
    end
    if (metaReset) begin
      r_resp_bits_taken <= 1'h0;
    end else if (io_resp_valid) begin
      r_resp_bits_taken <= io_resp_bits_taken;
    end
    if (metaReset) begin
      r_resp_bits_entry <= 5'h0;
    end else if (io_resp_valid) begin
      r_resp_bits_entry <= io_resp_bits_entry;
    end
    if (metaReset) begin
      _T_1163 <= 8'h0;
    end else if (io_bht_update_valid) begin
      if (io_bht_update_bits_branch) begin
        if (io_bht_update_bits_mispredict) begin
          _T_1163 <= _T_1247;
        end else if (io_bht_advance_valid) begin
          _T_1163 <= _T_1235;
        end
      end else if (io_bht_update_bits_mispredict) begin
        _T_1163 <= io_bht_update_bits_prediction_history;
      end else if (io_bht_advance_valid) begin
        _T_1163 <= _T_1235;
      end
    end else if (io_bht_advance_valid) begin
      _T_1163 <= _T_1235;
    end
    if (metaReset) begin
      _T_1252 <= 3'h0;
    end else if (io_ras_update_valid) begin
      if (_T_1331) begin
        if (_T_1332) begin
          _T_1252 <= _T_1334;
        end
      end else if (_T_1341) begin
        if (~_T_1324) begin
          _T_1252 <= _T_1346;
        end
      end
    end
    if (metaReset) begin
      _T_1254 <= 3'h0;
    end else if (io_ras_update_valid) begin
      if (_T_1331) begin
        if (_T_1335) begin
          _T_1254 <= _T_1338;
        end else begin
          _T_1254 <= 3'h0;
        end
      end else if (_T_1341) begin
        if (~_T_1324) begin
          if (_T_1347) begin
            _T_1254 <= _T_1351;
          end else begin
            _T_1254 <= 3'h5;
          end
        end
      end
    end
    if (metaReset) begin
      _T_1258_0 <= 39'h0;
    end else if (io_ras_update_valid) begin
      if (_T_1331) begin
        if (3'h0 == _T_1339) begin
          _T_1258_0 <= io_ras_update_bits_returnAddr;
        end
      end
    end
    if (metaReset) begin
      _T_1258_1 <= 39'h0;
    end else if (io_ras_update_valid) begin
      if (_T_1331) begin
        if (3'h1 == _T_1339) begin
          _T_1258_1 <= io_ras_update_bits_returnAddr;
        end
      end
    end
    if (metaReset) begin
      _T_1258_2 <= 39'h0;
    end else if (io_ras_update_valid) begin
      if (_T_1331) begin
        if (3'h2 == _T_1339) begin
          _T_1258_2 <= io_ras_update_bits_returnAddr;
        end
      end
    end
    if (metaReset) begin
      _T_1258_3 <= 39'h0;
    end else if (io_ras_update_valid) begin
      if (_T_1331) begin
        if (3'h3 == _T_1339) begin
          _T_1258_3 <= io_ras_update_bits_returnAddr;
        end
      end
    end
    if (metaReset) begin
      _T_1258_4 <= 39'h0;
    end else if (io_ras_update_valid) begin
      if (_T_1331) begin
        if (3'h4 == _T_1339) begin
          _T_1258_4 <= io_ras_update_bits_returnAddr;
        end
      end
    end
    if (metaReset) begin
      _T_1258_5 <= 39'h0;
    end else if (io_ras_update_valid) begin
      if (_T_1331) begin
        if (3'h5 == _T_1339) begin
          _T_1258_5 <= io_ras_update_bits_returnAddr;
        end
      end
    end
    BTB_state <= BTB_xor0;
    if (!(BTB_cov_read_data)) begin
      BTB_covSum <= BTB_covSum + 1'h1;
    end
  end
  always @(posedge clock) begin
    if(BTB_cov_write_en & BTB_cov_write_mask) begin
      BTB_cov[BTB_cov_write_addr] <= BTB_cov_write_data; // @[Coverage map for BTB]
    end
  end
endmodule
module TLMonitor_66(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_param,
  input  [3:0]  io_in_a_bits_size,
  input  [1:0]  io_in_a_bits_source,
  input  [31:0] io_in_a_bits_address,
  input  [7:0]  io_in_a_bits_mask,
  input         io_in_a_bits_corrupt,
  input         io_in_b_ready,
  input         io_in_b_valid,
  input  [2:0]  io_in_b_bits_opcode,
  input  [1:0]  io_in_b_bits_param,
  input  [3:0]  io_in_b_bits_size,
  input  [1:0]  io_in_b_bits_source,
  input  [31:0] io_in_b_bits_address,
  input  [7:0]  io_in_b_bits_mask,
  input         io_in_b_bits_corrupt,
  input         io_in_c_ready,
  input         io_in_c_valid,
  input  [2:0]  io_in_c_bits_opcode,
  input  [2:0]  io_in_c_bits_param,
  input  [3:0]  io_in_c_bits_size,
  input  [1:0]  io_in_c_bits_source,
  input  [31:0] io_in_c_bits_address,
  input         io_in_d_ready,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [1:0]  io_in_d_bits_param,
  input  [3:0]  io_in_d_bits_size,
  input  [1:0]  io_in_d_bits_source,
  input  [1:0]  io_in_d_bits_sink,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt,
  input         io_in_e_ready,
  input         io_in_e_valid,
  input  [1:0]  io_in_e_bits_sink,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire  _T_20; // @[Parameters.scala 44:9]
  wire  _T_21; // @[Parameters.scala 44:9]
  wire  _T_22; // @[Parameters.scala 44:9]
  wire  _T_32; // @[Parameters.scala 280:46]
  wire  _T_33; // @[Parameters.scala 280:46]
  wire [26:0] _T_35; // @[package.scala 185:77]
  wire [31:0] _GEN_33; // @[Edges.scala 21:16]
  wire [31:0] _T_38; // @[Edges.scala 21:16]
  wire  _T_39; // @[Edges.scala 21:24]
  wire [3:0] _T_42; // @[OneHot.scala 52:12]
  wire [2:0] _T_44; // @[Misc.scala 206:81]
  wire  _T_45; // @[Misc.scala 210:21]
  wire  _T_50; // @[Misc.scala 219:38]
  wire  _T_51; // @[Misc.scala 219:29]
  wire  _T_53; // @[Misc.scala 219:38]
  wire  _T_54; // @[Misc.scala 219:29]
  wire  _T_58; // @[Misc.scala 218:27]
  wire  _T_59; // @[Misc.scala 219:38]
  wire  _T_60; // @[Misc.scala 219:29]
  wire  _T_61; // @[Misc.scala 218:27]
  wire  _T_62; // @[Misc.scala 219:38]
  wire  _T_63; // @[Misc.scala 219:29]
  wire  _T_64; // @[Misc.scala 218:27]
  wire  _T_65; // @[Misc.scala 219:38]
  wire  _T_66; // @[Misc.scala 219:29]
  wire  _T_67; // @[Misc.scala 218:27]
  wire  _T_68; // @[Misc.scala 219:38]
  wire  _T_69; // @[Misc.scala 219:29]
  wire  _T_73; // @[Misc.scala 218:27]
  wire  _T_74; // @[Misc.scala 219:38]
  wire  _T_75; // @[Misc.scala 219:29]
  wire  _T_76; // @[Misc.scala 218:27]
  wire  _T_77; // @[Misc.scala 219:38]
  wire  _T_78; // @[Misc.scala 219:29]
  wire  _T_79; // @[Misc.scala 218:27]
  wire  _T_80; // @[Misc.scala 219:38]
  wire  _T_81; // @[Misc.scala 219:29]
  wire  _T_82; // @[Misc.scala 218:27]
  wire  _T_83; // @[Misc.scala 219:38]
  wire  _T_84; // @[Misc.scala 219:29]
  wire  _T_85; // @[Misc.scala 218:27]
  wire  _T_86; // @[Misc.scala 219:38]
  wire  _T_87; // @[Misc.scala 219:29]
  wire  _T_88; // @[Misc.scala 218:27]
  wire  _T_89; // @[Misc.scala 219:38]
  wire  _T_90; // @[Misc.scala 219:29]
  wire  _T_91; // @[Misc.scala 218:27]
  wire  _T_92; // @[Misc.scala 219:38]
  wire  _T_93; // @[Misc.scala 219:29]
  wire  _T_94; // @[Misc.scala 218:27]
  wire  _T_95; // @[Misc.scala 219:38]
  wire  _T_96; // @[Misc.scala 219:29]
  wire [7:0] _T_103; // @[Cat.scala 30:58]
  wire [32:0] _T_107; // @[Parameters.scala 121:49]
  wire  _T_133; // @[Monitor.scala 48:25]
  wire  _T_135; // @[Parameters.scala 90:42]
  wire [31:0] _T_138; // @[Parameters.scala 121:31]
  wire [32:0] _T_139; // @[Parameters.scala 121:49]
  wire [32:0] _T_141; // @[Parameters.scala 121:52]
  wire  _T_142; // @[Parameters.scala 121:67]
  wire  _T_143; // @[Parameters.scala 168:56]
  wire [31:0] _T_145; // @[Parameters.scala 121:31]
  wire [32:0] _T_146; // @[Parameters.scala 121:49]
  wire [32:0] _T_148; // @[Parameters.scala 121:52]
  wire  _T_149; // @[Parameters.scala 121:67]
  wire [31:0] _T_150; // @[Parameters.scala 121:31]
  wire [32:0] _T_151; // @[Parameters.scala 121:49]
  wire [32:0] _T_153; // @[Parameters.scala 121:52]
  wire  _T_154; // @[Parameters.scala 121:67]
  wire [31:0] _T_155; // @[Parameters.scala 121:31]
  wire [32:0] _T_156; // @[Parameters.scala 121:49]
  wire [32:0] _T_158; // @[Parameters.scala 121:52]
  wire  _T_159; // @[Parameters.scala 121:67]
  wire [32:0] _T_163; // @[Parameters.scala 121:52]
  wire  _T_164; // @[Parameters.scala 121:67]
  wire [31:0] _T_165; // @[Parameters.scala 121:31]
  wire [32:0] _T_166; // @[Parameters.scala 121:49]
  wire [32:0] _T_168; // @[Parameters.scala 121:52]
  wire  _T_169; // @[Parameters.scala 121:67]
  wire [31:0] _T_170; // @[Parameters.scala 121:31]
  wire [32:0] _T_171; // @[Parameters.scala 121:49]
  wire [32:0] _T_173; // @[Parameters.scala 121:52]
  wire  _T_174; // @[Parameters.scala 121:67]
  wire  _T_175; // @[Parameters.scala 169:42]
  wire  _T_176; // @[Parameters.scala 169:42]
  wire  _T_177; // @[Parameters.scala 169:42]
  wire  _T_184; // @[Monitor.scala 49:14]
  wire  _T_198; // @[Parameters.scala 89:48]
  wire  _T_200; // @[Mux.scala 19:72]
  wire  _T_208; // @[Monitor.scala 50:14]
  wire  _T_211; // @[Monitor.scala 51:14]
  wire  _T_215; // @[Monitor.scala 52:14]
  wire  _T_218; // @[Monitor.scala 53:14]
  wire  _T_220; // @[Bundles.scala 109:27]
  wire  _T_222; // @[Monitor.scala 54:14]
  wire  _T_225; // @[Monitor.scala 55:28]
  wire  _T_227; // @[Monitor.scala 55:14]
  wire  _T_231; // @[Monitor.scala 56:14]
  wire  _T_233; // @[Monitor.scala 59:25]
  wire  _T_324; // @[Monitor.scala 66:28]
  wire  _T_326; // @[Monitor.scala 66:14]
  wire  _T_337; // @[Monitor.scala 71:25]
  wire  _T_339; // @[Parameters.scala 90:42]
  wire  _T_347; // @[Parameters.scala 168:56]
  wire  _T_382; // @[Parameters.scala 169:42]
  wire  _T_383; // @[Parameters.scala 169:42]
  wire  _T_384; // @[Parameters.scala 169:42]
  wire  _T_385; // @[Parameters.scala 169:42]
  wire  _T_386; // @[Parameters.scala 169:42]
  wire  _T_387; // @[Parameters.scala 168:56]
  wire  _T_389; // @[Parameters.scala 170:30]
  wire  _T_391; // @[Monitor.scala 72:14]
  wire  _T_399; // @[Monitor.scala 75:28]
  wire  _T_401; // @[Monitor.scala 75:14]
  wire  _T_403; // @[Monitor.scala 76:27]
  wire  _T_405; // @[Monitor.scala 76:14]
  wire  _T_411; // @[Monitor.scala 80:25]
  wire  _T_448; // @[Parameters.scala 169:42]
  wire  _T_449; // @[Parameters.scala 168:56]
  wire  _T_451; // @[Parameters.scala 90:42]
  wire  _T_459; // @[Parameters.scala 168:56]
  wire  _T_468; // @[Parameters.scala 170:30]
  wire  _T_469; // @[Parameters.scala 170:30]
  wire  _T_472; // @[Monitor.scala 81:14]
  wire  _T_488; // @[Monitor.scala 88:25]
  wire [7:0] _T_562; // @[Monitor.scala 93:28]
  wire  _T_563; // @[Monitor.scala 93:37]
  wire  _T_565; // @[Monitor.scala 93:14]
  wire  _T_567; // @[Monitor.scala 96:25]
  wire  _T_569; // @[Parameters.scala 90:42]
  wire  _T_595; // @[Parameters.scala 168:56]
  wire  _T_618; // @[Monitor.scala 97:14]
  wire  _T_626; // @[Bundles.scala 139:33]
  wire  _T_628; // @[Monitor.scala 100:14]
  wire  _T_634; // @[Monitor.scala 104:25]
  wire  _T_693; // @[Bundles.scala 146:30]
  wire  _T_695; // @[Monitor.scala 108:14]
  wire  _T_701; // @[Monitor.scala 112:25]
  wire  _T_752; // @[Monitor.scala 113:14]
  wire  _T_768; // @[Bundles.scala 43:24]
  wire  _T_770; // @[Monitor.scala 268:12]
  wire  _T_772; // @[Parameters.scala 44:9]
  wire  _T_773; // @[Parameters.scala 44:9]
  wire  _T_774; // @[Parameters.scala 44:9]
  wire  _T_784; // @[Parameters.scala 280:46]
  wire  _T_785; // @[Parameters.scala 280:46]
  wire  _T_787; // @[Monitor.scala 275:25]
  wire  _T_789; // @[Monitor.scala 276:14]
  wire  _T_791; // @[Monitor.scala 277:27]
  wire  _T_793; // @[Monitor.scala 277:14]
  wire  _T_795; // @[Monitor.scala 278:28]
  wire  _T_797; // @[Monitor.scala 278:14]
  wire  _T_801; // @[Monitor.scala 279:14]
  wire  _T_805; // @[Monitor.scala 280:14]
  wire  _T_807; // @[Monitor.scala 283:25]
  wire  _T_818; // @[Bundles.scala 103:26]
  wire  _T_820; // @[Monitor.scala 287:14]
  wire  _T_822; // @[Monitor.scala 288:28]
  wire  _T_824; // @[Monitor.scala 288:14]
  wire  _T_835; // @[Monitor.scala 293:25]
  wire  _T_855; // @[Monitor.scala 299:30]
  wire  _T_857; // @[Monitor.scala 299:14]
  wire  _T_864; // @[Monitor.scala 303:25]
  wire  _T_881; // @[Monitor.scala 311:25]
  wire  _T_899; // @[Monitor.scala 319:25]
  wire  _T_916; // @[Bundles.scala 41:24]
  wire  _T_918; // @[Monitor.scala 122:12]
  wire  _T_920; // @[Parameters.scala 44:9]
  wire [32:0] _T_923; // @[Parameters.scala 121:49]
  wire  _T_928; // @[Parameters.scala 44:9]
  wire  _T_936; // @[Parameters.scala 44:9]
  wire [31:0] _T_949; // @[Parameters.scala 121:31]
  wire [32:0] _T_950; // @[Parameters.scala 121:49]
  wire [32:0] _T_952; // @[Parameters.scala 121:52]
  wire  _T_953; // @[Parameters.scala 121:67]
  wire [31:0] _T_954; // @[Parameters.scala 121:31]
  wire [32:0] _T_955; // @[Parameters.scala 121:49]
  wire [32:0] _T_957; // @[Parameters.scala 121:52]
  wire  _T_958; // @[Parameters.scala 121:67]
  wire [31:0] _T_959; // @[Parameters.scala 121:31]
  wire [32:0] _T_960; // @[Parameters.scala 121:49]
  wire [32:0] _T_962; // @[Parameters.scala 121:52]
  wire  _T_963; // @[Parameters.scala 121:67]
  wire [32:0] _T_967; // @[Parameters.scala 121:52]
  wire  _T_968; // @[Parameters.scala 121:67]
  wire [31:0] _T_969; // @[Parameters.scala 121:31]
  wire [32:0] _T_970; // @[Parameters.scala 121:49]
  wire [32:0] _T_972; // @[Parameters.scala 121:52]
  wire  _T_973; // @[Parameters.scala 121:67]
  wire [31:0] _T_974; // @[Parameters.scala 121:31]
  wire [32:0] _T_975; // @[Parameters.scala 121:49]
  wire [32:0] _T_977; // @[Parameters.scala 121:52]
  wire  _T_978; // @[Parameters.scala 121:67]
  wire [31:0] _T_979; // @[Parameters.scala 121:31]
  wire [32:0] _T_980; // @[Parameters.scala 121:49]
  wire [32:0] _T_982; // @[Parameters.scala 121:52]
  wire  _T_983; // @[Parameters.scala 121:67]
  wire  _T_997; // @[Parameters.scala 155:64]
  wire  _T_998; // @[Parameters.scala 155:64]
  wire  _T_999; // @[Parameters.scala 155:64]
  wire  _T_1000; // @[Parameters.scala 155:64]
  wire  _T_1001; // @[Parameters.scala 155:64]
  wire  _T_1002; // @[Parameters.scala 155:64]
  wire [26:0] _T_1004; // @[package.scala 185:77]
  wire [31:0] _GEN_34; // @[Edges.scala 21:16]
  wire [31:0] _T_1007; // @[Edges.scala 21:16]
  wire  _T_1008; // @[Edges.scala 21:24]
  wire [3:0] _T_1011; // @[OneHot.scala 52:12]
  wire [2:0] _T_1013; // @[Misc.scala 206:81]
  wire  _T_1014; // @[Misc.scala 210:21]
  wire  _T_1019; // @[Misc.scala 219:38]
  wire  _T_1020; // @[Misc.scala 219:29]
  wire  _T_1022; // @[Misc.scala 219:38]
  wire  _T_1023; // @[Misc.scala 219:29]
  wire  _T_1027; // @[Misc.scala 218:27]
  wire  _T_1028; // @[Misc.scala 219:38]
  wire  _T_1029; // @[Misc.scala 219:29]
  wire  _T_1030; // @[Misc.scala 218:27]
  wire  _T_1031; // @[Misc.scala 219:38]
  wire  _T_1032; // @[Misc.scala 219:29]
  wire  _T_1033; // @[Misc.scala 218:27]
  wire  _T_1034; // @[Misc.scala 219:38]
  wire  _T_1035; // @[Misc.scala 219:29]
  wire  _T_1036; // @[Misc.scala 218:27]
  wire  _T_1037; // @[Misc.scala 219:38]
  wire  _T_1038; // @[Misc.scala 219:29]
  wire  _T_1042; // @[Misc.scala 218:27]
  wire  _T_1043; // @[Misc.scala 219:38]
  wire  _T_1044; // @[Misc.scala 219:29]
  wire  _T_1045; // @[Misc.scala 218:27]
  wire  _T_1046; // @[Misc.scala 219:38]
  wire  _T_1047; // @[Misc.scala 219:29]
  wire  _T_1048; // @[Misc.scala 218:27]
  wire  _T_1049; // @[Misc.scala 219:38]
  wire  _T_1050; // @[Misc.scala 219:29]
  wire  _T_1051; // @[Misc.scala 218:27]
  wire  _T_1052; // @[Misc.scala 219:38]
  wire  _T_1053; // @[Misc.scala 219:29]
  wire  _T_1054; // @[Misc.scala 218:27]
  wire  _T_1055; // @[Misc.scala 219:38]
  wire  _T_1056; // @[Misc.scala 219:29]
  wire  _T_1057; // @[Misc.scala 218:27]
  wire  _T_1058; // @[Misc.scala 219:38]
  wire  _T_1059; // @[Misc.scala 219:29]
  wire  _T_1060; // @[Misc.scala 218:27]
  wire  _T_1061; // @[Misc.scala 219:38]
  wire  _T_1062; // @[Misc.scala 219:29]
  wire  _T_1063; // @[Misc.scala 218:27]
  wire  _T_1064; // @[Misc.scala 219:38]
  wire  _T_1065; // @[Misc.scala 219:29]
  wire [7:0] _T_1072; // @[Cat.scala 30:58]
  wire [1:0] _T_1088; // @[Mux.scala 19:72]
  wire [1:0] _GEN_35; // @[Mux.scala 19:72]
  wire [1:0] _T_1090; // @[Mux.scala 19:72]
  wire  _T_1093; // @[Monitor.scala 130:117]
  wire  _T_1094; // @[Monitor.scala 132:25]
  wire  _T_1107; // @[Parameters.scala 89:48]
  wire  _T_1109; // @[Mux.scala 19:72]
  wire  _T_1117; // @[Monitor.scala 133:14]
  wire  _T_1120; // @[Monitor.scala 134:14]
  wire  _T_1123; // @[Monitor.scala 135:14]
  wire  _T_1126; // @[Monitor.scala 136:14]
  wire  _T_1128; // @[Bundles.scala 103:26]
  wire  _T_1130; // @[Monitor.scala 137:14]
  wire  _T_1132; // @[Monitor.scala 138:27]
  wire  _T_1134; // @[Monitor.scala 138:14]
  wire  _T_1138; // @[Monitor.scala 139:14]
  wire  _T_1140; // @[Monitor.scala 142:25]
  wire  _T_1153; // @[Monitor.scala 147:28]
  wire  _T_1155; // @[Monitor.scala 147:14]
  wire  _T_1165; // @[Monitor.scala 152:25]
  wire  _T_1186; // @[Monitor.scala 161:25]
  wire [7:0] _T_1204; // @[Monitor.scala 167:28]
  wire  _T_1205; // @[Monitor.scala 167:37]
  wire  _T_1207; // @[Monitor.scala 167:14]
  wire  _T_1209; // @[Monitor.scala 170:25]
  wire  _T_1230; // @[Monitor.scala 179:25]
  wire  _T_1251; // @[Monitor.scala 188:25]
  wire  _T_1276; // @[Parameters.scala 44:9]
  wire  _T_1277; // @[Parameters.scala 44:9]
  wire  _T_1278; // @[Parameters.scala 44:9]
  wire  _T_1288; // @[Parameters.scala 280:46]
  wire  _T_1289; // @[Parameters.scala 280:46]
  wire [26:0] _T_1291; // @[package.scala 185:77]
  wire [31:0] _GEN_36; // @[Edges.scala 21:16]
  wire [31:0] _T_1294; // @[Edges.scala 21:16]
  wire  _T_1295; // @[Edges.scala 21:24]
  wire [31:0] _T_1296; // @[Parameters.scala 121:31]
  wire [32:0] _T_1297; // @[Parameters.scala 121:49]
  wire [32:0] _T_1299; // @[Parameters.scala 121:52]
  wire  _T_1300; // @[Parameters.scala 121:67]
  wire [31:0] _T_1301; // @[Parameters.scala 121:31]
  wire [32:0] _T_1302; // @[Parameters.scala 121:49]
  wire [32:0] _T_1304; // @[Parameters.scala 121:52]
  wire  _T_1305; // @[Parameters.scala 121:67]
  wire [31:0] _T_1306; // @[Parameters.scala 121:31]
  wire [32:0] _T_1307; // @[Parameters.scala 121:49]
  wire [32:0] _T_1309; // @[Parameters.scala 121:52]
  wire  _T_1310; // @[Parameters.scala 121:67]
  wire [32:0] _T_1312; // @[Parameters.scala 121:49]
  wire [32:0] _T_1314; // @[Parameters.scala 121:52]
  wire  _T_1315; // @[Parameters.scala 121:67]
  wire [31:0] _T_1316; // @[Parameters.scala 121:31]
  wire [32:0] _T_1317; // @[Parameters.scala 121:49]
  wire [32:0] _T_1319; // @[Parameters.scala 121:52]
  wire  _T_1320; // @[Parameters.scala 121:67]
  wire [31:0] _T_1321; // @[Parameters.scala 121:31]
  wire [32:0] _T_1322; // @[Parameters.scala 121:49]
  wire [32:0] _T_1324; // @[Parameters.scala 121:52]
  wire  _T_1325; // @[Parameters.scala 121:67]
  wire [31:0] _T_1326; // @[Parameters.scala 121:31]
  wire [32:0] _T_1327; // @[Parameters.scala 121:49]
  wire [32:0] _T_1329; // @[Parameters.scala 121:52]
  wire  _T_1330; // @[Parameters.scala 121:67]
  wire  _T_1344; // @[Parameters.scala 155:64]
  wire  _T_1345; // @[Parameters.scala 155:64]
  wire  _T_1346; // @[Parameters.scala 155:64]
  wire  _T_1347; // @[Parameters.scala 155:64]
  wire  _T_1348; // @[Parameters.scala 155:64]
  wire  _T_1349; // @[Parameters.scala 155:64]
  wire  _T_1379; // @[Monitor.scala 207:25]
  wire  _T_1381; // @[Monitor.scala 208:14]
  wire  _T_1384; // @[Monitor.scala 209:14]
  wire  _T_1386; // @[Monitor.scala 210:27]
  wire  _T_1388; // @[Monitor.scala 210:14]
  wire  _T_1391; // @[Monitor.scala 211:14]
  wire  _T_1393; // @[Bundles.scala 121:29]
  wire  _T_1395; // @[Monitor.scala 212:14]
  wire  _T_1401; // @[Monitor.scala 216:25]
  wire  _T_1419; // @[Monitor.scala 224:25]
  wire  _T_1421; // @[Parameters.scala 90:42]
  wire  _T_1429; // @[Parameters.scala 168:56]
  wire  _T_1470; // @[Monitor.scala 225:14]
  wire  _T_1484; // @[Parameters.scala 89:48]
  wire  _T_1486; // @[Mux.scala 19:72]
  wire  _T_1494; // @[Monitor.scala 226:14]
  wire  _T_1506; // @[Bundles.scala 115:29]
  wire  _T_1508; // @[Monitor.scala 230:14]
  wire  _T_1514; // @[Monitor.scala 234:25]
  wire  _T_1605; // @[Monitor.scala 243:25]
  wire  _T_1615; // @[Monitor.scala 247:28]
  wire  _T_1617; // @[Monitor.scala 247:14]
  wire  _T_1623; // @[Monitor.scala 251:25]
  wire  _T_1637; // @[Monitor.scala 258:25]
  wire  _T_1659; // @[Bundles.scala 277:22]
  wire [8:0] _T_1664; // @[Edges.scala 220:59]
  reg [8:0] _T_1669; // @[Edges.scala 229:27]
  reg [31:0] _RAND_0;
  wire [8:0] _T_1672; // @[Edges.scala 230:28]
  wire  _T_1673; // @[Edges.scala 231:25]
  reg [2:0] _T_1682; // @[Monitor.scala 349:22]
  reg [31:0] _RAND_1;
  reg [2:0] _T_1684; // @[Monitor.scala 350:22]
  reg [31:0] _RAND_2;
  reg [3:0] _T_1686; // @[Monitor.scala 351:22]
  reg [31:0] _RAND_3;
  reg [1:0] _T_1688; // @[Monitor.scala 352:22]
  reg [31:0] _RAND_4;
  reg [31:0] _T_1690; // @[Monitor.scala 353:22]
  reg [31:0] _RAND_5;
  wire  _T_1692; // @[Monitor.scala 354:19]
  wire  _T_1693; // @[Monitor.scala 355:29]
  wire  _T_1695; // @[Monitor.scala 355:14]
  wire  _T_1697; // @[Monitor.scala 356:29]
  wire  _T_1699; // @[Monitor.scala 356:14]
  wire  _T_1701; // @[Monitor.scala 357:29]
  wire  _T_1703; // @[Monitor.scala 357:14]
  wire  _T_1705; // @[Monitor.scala 358:29]
  wire  _T_1707; // @[Monitor.scala 358:14]
  wire  _T_1709; // @[Monitor.scala 359:29]
  wire  _T_1711; // @[Monitor.scala 359:14]
  wire  _T_1714; // @[Monitor.scala 361:20]
  wire  _T_1715; // @[Bundles.scala 277:22]
  wire [26:0] _T_1717; // @[package.scala 185:77]
  wire [8:0] _T_1720; // @[Edges.scala 220:59]
  reg [8:0] _T_1724; // @[Edges.scala 229:27]
  reg [31:0] _RAND_6;
  wire [8:0] _T_1727; // @[Edges.scala 230:28]
  wire  _T_1728; // @[Edges.scala 231:25]
  reg [2:0] _T_1737; // @[Monitor.scala 418:22]
  reg [31:0] _RAND_7;
  reg [1:0] _T_1739; // @[Monitor.scala 419:22]
  reg [31:0] _RAND_8;
  reg [3:0] _T_1741; // @[Monitor.scala 420:22]
  reg [31:0] _RAND_9;
  reg [1:0] _T_1743; // @[Monitor.scala 421:22]
  reg [31:0] _RAND_10;
  reg [1:0] _T_1745; // @[Monitor.scala 422:22]
  reg [31:0] _RAND_11;
  reg  _T_1747; // @[Monitor.scala 423:22]
  reg [31:0] _RAND_12;
  wire  _T_1749; // @[Monitor.scala 424:19]
  wire  _T_1750; // @[Monitor.scala 425:29]
  wire  _T_1752; // @[Monitor.scala 425:14]
  wire  _T_1754; // @[Monitor.scala 426:29]
  wire  _T_1756; // @[Monitor.scala 426:14]
  wire  _T_1758; // @[Monitor.scala 427:29]
  wire  _T_1760; // @[Monitor.scala 427:14]
  wire  _T_1762; // @[Monitor.scala 428:29]
  wire  _T_1764; // @[Monitor.scala 428:14]
  wire  _T_1766; // @[Monitor.scala 429:29]
  wire  _T_1768; // @[Monitor.scala 429:14]
  wire  _T_1770; // @[Monitor.scala 430:29]
  wire  _T_1772; // @[Monitor.scala 430:14]
  wire  _T_1775; // @[Monitor.scala 432:20]
  wire  _T_1776; // @[Bundles.scala 277:22]
  reg [8:0] _T_1786; // @[Edges.scala 229:27]
  reg [31:0] _RAND_13;
  wire [8:0] _T_1789; // @[Edges.scala 230:28]
  wire  _T_1790; // @[Edges.scala 231:25]
  reg [2:0] _T_1799; // @[Monitor.scala 372:22]
  reg [31:0] _RAND_14;
  reg [1:0] _T_1801; // @[Monitor.scala 373:22]
  reg [31:0] _RAND_15;
  reg [3:0] _T_1803; // @[Monitor.scala 374:22]
  reg [31:0] _RAND_16;
  reg [1:0] _T_1805; // @[Monitor.scala 375:22]
  reg [31:0] _RAND_17;
  reg [31:0] _T_1807; // @[Monitor.scala 376:22]
  reg [31:0] _RAND_18;
  wire  _T_1809; // @[Monitor.scala 377:19]
  wire  _T_1810; // @[Monitor.scala 378:29]
  wire  _T_1812; // @[Monitor.scala 378:14]
  wire  _T_1814; // @[Monitor.scala 379:29]
  wire  _T_1816; // @[Monitor.scala 379:14]
  wire  _T_1818; // @[Monitor.scala 380:29]
  wire  _T_1820; // @[Monitor.scala 380:14]
  wire  _T_1822; // @[Monitor.scala 381:29]
  wire  _T_1824; // @[Monitor.scala 381:14]
  wire  _T_1826; // @[Monitor.scala 382:29]
  wire  _T_1828; // @[Monitor.scala 382:14]
  wire  _T_1831; // @[Monitor.scala 384:20]
  wire  _T_1832; // @[Bundles.scala 277:22]
  wire [8:0] _T_1837; // @[Edges.scala 220:59]
  reg [8:0] _T_1841; // @[Edges.scala 229:27]
  reg [31:0] _RAND_19;
  wire [8:0] _T_1844; // @[Edges.scala 230:28]
  wire  _T_1845; // @[Edges.scala 231:25]
  reg [2:0] _T_1854; // @[Monitor.scala 395:22]
  reg [31:0] _RAND_20;
  reg [2:0] _T_1856; // @[Monitor.scala 396:22]
  reg [31:0] _RAND_21;
  reg [3:0] _T_1858; // @[Monitor.scala 397:22]
  reg [31:0] _RAND_22;
  reg [1:0] _T_1860; // @[Monitor.scala 398:22]
  reg [31:0] _RAND_23;
  reg [31:0] _T_1862; // @[Monitor.scala 399:22]
  reg [31:0] _RAND_24;
  wire  _T_1864; // @[Monitor.scala 400:19]
  wire  _T_1865; // @[Monitor.scala 401:29]
  wire  _T_1867; // @[Monitor.scala 401:14]
  wire  _T_1869; // @[Monitor.scala 402:29]
  wire  _T_1871; // @[Monitor.scala 402:14]
  wire  _T_1873; // @[Monitor.scala 403:29]
  wire  _T_1875; // @[Monitor.scala 403:14]
  wire  _T_1877; // @[Monitor.scala 404:29]
  wire  _T_1879; // @[Monitor.scala 404:14]
  wire  _T_1881; // @[Monitor.scala 405:29]
  wire  _T_1883; // @[Monitor.scala 405:14]
  wire  _T_1886; // @[Monitor.scala 407:20]
  reg [2:0] _T_1888; // @[Monitor.scala 452:27]
  reg [31:0] _RAND_25;
  reg [8:0] _T_1899; // @[Edges.scala 229:27]
  reg [31:0] _RAND_26;
  wire [8:0] _T_1902; // @[Edges.scala 230:28]
  wire  _T_1903; // @[Edges.scala 231:25]
  reg [8:0] _T_1920; // @[Edges.scala 229:27]
  reg [31:0] _RAND_27;
  wire [8:0] _T_1923; // @[Edges.scala 230:28]
  wire  _T_1924; // @[Edges.scala 231:25]
  wire  _T_1935; // @[Monitor.scala 458:27]
  wire [3:0] _T_1937; // @[OneHot.scala 45:35]
  wire [2:0] _T_1938; // @[Monitor.scala 460:23]
  wire  _T_1942; // @[Monitor.scala 460:13]
  wire [3:0] _GEN_27; // @[Monitor.scala 458:72]
  wire  _T_1948; // @[Monitor.scala 465:27]
  wire  _T_1951; // @[Monitor.scala 465:72]
  wire [3:0] _T_1952; // @[OneHot.scala 45:35]
  wire [2:0] _T_1953; // @[Monitor.scala 467:21]
  wire [2:0] _T_1954; // @[Monitor.scala 467:32]
  wire  _T_1957; // @[Monitor.scala 467:13]
  wire [3:0] _GEN_28; // @[Monitor.scala 465:91]
  wire  _T_1959; // @[Monitor.scala 471:20]
  wire  _T_1960; // @[Monitor.scala 471:40]
  wire  _T_1962; // @[Monitor.scala 471:30]
  wire  _T_1964; // @[Monitor.scala 471:13]
  wire [2:0] _T_1966; // @[Monitor.scala 474:27]
  wire [2:0] _T_1968; // @[Monitor.scala 474:36]
  reg [3:0] _T_1986; // @[Monitor.scala 486:27]
  reg [31:0] _RAND_28;
  reg [8:0] _T_1996; // @[Edges.scala 229:27]
  reg [31:0] _RAND_29;
  wire [8:0] _T_1999; // @[Edges.scala 230:28]
  wire  _T_2000; // @[Edges.scala 231:25]
  wire  _T_2011; // @[Monitor.scala 492:27]
  wire  _T_2015; // @[Edges.scala 71:40]
  wire  _T_2016; // @[Monitor.scala 492:38]
  wire [3:0] _T_2017; // @[OneHot.scala 45:35]
  wire [3:0] _T_2018; // @[Monitor.scala 494:23]
  wire  _T_2022; // @[Monitor.scala 494:13]
  wire [3:0] _GEN_31; // @[Monitor.scala 492:72]
  wire  _T_2026; // @[Bundles.scala 277:22]
  wire [3:0] _T_2029; // @[OneHot.scala 45:35]
  wire [3:0] _T_2030; // @[Monitor.scala 500:21]
  wire [3:0] _T_2031; // @[Monitor.scala 500:32]
  wire  _T_2034; // @[Monitor.scala 500:13]
  wire [3:0] _GEN_32; // @[Monitor.scala 498:73]
  wire [3:0] _T_2036; // @[Monitor.scala 505:27]
  wire [3:0] _T_2038; // @[Monitor.scala 505:36]
  wire  _GEN_37; // @[Monitor.scala 49:14]
  wire  _GEN_53; // @[Monitor.scala 60:14]
  wire  _GEN_71; // @[Monitor.scala 72:14]
  wire  _GEN_83; // @[Monitor.scala 81:14]
  wire  _GEN_93; // @[Monitor.scala 89:14]
  wire  _GEN_103; // @[Monitor.scala 97:14]
  wire  _GEN_113; // @[Monitor.scala 105:14]
  wire  _GEN_123; // @[Monitor.scala 113:14]
  wire  _GEN_133; // @[Monitor.scala 276:14]
  wire  _GEN_143; // @[Monitor.scala 284:14]
  wire  _GEN_153; // @[Monitor.scala 294:14]
  wire  _GEN_163; // @[Monitor.scala 304:14]
  wire  _GEN_169; // @[Monitor.scala 312:14]
  wire  _GEN_175; // @[Monitor.scala 320:14]
  wire  _GEN_181; // @[Monitor.scala 133:14]
  wire  _GEN_195; // @[Monitor.scala 143:14]
  wire  _GEN_209; // @[Monitor.scala 153:14]
  wire  _GEN_221; // @[Monitor.scala 162:14]
  wire  _GEN_233; // @[Monitor.scala 171:14]
  wire  _GEN_243; // @[Monitor.scala 180:14]
  wire  _GEN_253; // @[Monitor.scala 189:14]
  wire  _GEN_265; // @[Monitor.scala 208:14]
  wire  _GEN_275; // @[Monitor.scala 217:14]
  wire  _GEN_285; // @[Monitor.scala 225:14]
  wire  _GEN_297; // @[Monitor.scala 235:14]
  wire  _GEN_309; // @[Monitor.scala 244:14]
  wire  _GEN_317; // @[Monitor.scala 252:14]
  wire  _GEN_325; // @[Monitor.scala 259:14]
  wire [29:0] TLMonitor_66_covSum;
  wire  stopEn0;
  wire  stopEn1;
  wire  stopEn2;
  wire  stopEn3;
  wire  stopEn4;
  wire  stopEn5;
  wire  stopEn6;
  wire  stopEn7;
  wire  stopEn8;
  wire  stopEn9;
  wire  stopEn10;
  wire  stopEn11;
  wire  stopEn12;
  wire  stopEn13;
  wire  stopEn14;
  wire  stopEn15;
  wire  stopEn16;
  wire  stopEn17;
  wire  stopEn18;
  wire  stopEn19;
  wire  stopEn20;
  wire  stopEn21;
  wire  stopEn22;
  wire  stopEn23;
  wire  stopEn24;
  wire  stopEn25;
  wire  stopEn26;
  wire  stopEn27;
  wire  stopEn28;
  wire  stopEn29;
  wire  stopEn30;
  wire  stopEn31;
  wire  stopEn32;
  wire  stopEn33;
  wire  stopEn34;
  wire  stopEn35;
  wire  stopEn36;
  wire  stopEn37;
  wire  stopEn38;
  wire  stopEn39;
  wire  stopEn40;
  wire  stopEn41;
  wire  stopEn42;
  wire  stopEn43;
  wire  stopEn44;
  wire  stopEn45;
  wire  stopEn46;
  wire  stopEn47;
  wire  stopEn48;
  wire  stopEn49;
  wire  stopEn50;
  wire  stopEn51;
  wire  stopEn52;
  wire  stopEn53;
  wire  stopEn54;
  wire  stopEn55;
  wire  stopEn56;
  wire  stopEn57;
  wire  stopEn58;
  wire  stopEn59;
  wire  stopEn60;
  wire  stopEn61;
  wire  stopEn62;
  wire  stopEn63;
  wire  stopEn64;
  wire  stopEn65;
  wire  stopEn66;
  wire  stopEn67;
  wire  stopEn68;
  wire  stopEn69;
  wire  stopEn70;
  wire  stopEn71;
  wire  stopEn72;
  wire  stopEn73;
  wire  stopEn74;
  wire  stopEn75;
  wire  stopEn76;
  wire  stopEn77;
  wire  stopEn78;
  wire  stopEn79;
  wire  stopEn80;
  wire  stopEn81;
  wire  stopEn82;
  wire  stopEn83;
  wire  stopEn84;
  wire  stopEn85;
  wire  stopEn86;
  wire  stopEn87;
  wire  stopEn88;
  wire  stopEn89;
  wire  stopEn90;
  wire  stopEn91;
  wire  stopEn92;
  wire  stopEn93;
  wire  stopEn94;
  wire  stopEn95;
  wire  stopEn96;
  wire  stopEn97;
  wire  stopEn98;
  wire  stopEn99;
  wire  stopEn100;
  wire  stopEn101;
  wire  stopEn102;
  wire  stopEn103;
  wire  stopEn104;
  wire  stopEn105;
  wire  stopEn106;
  wire  stopEn107;
  wire  stopEn108;
  wire  stopEn109;
  wire  stopEn110;
  wire  stopEn111;
  wire  stopEn112;
  wire  stopEn113;
  wire  stopEn114;
  wire  stopEn115;
  wire  stopEn116;
  wire  stopEn117;
  wire  stopEn118;
  wire  stopEn119;
  wire  stopEn120;
  wire  stopEn121;
  wire  stopEn122;
  wire  stopEn123;
  wire  stopEn124;
  wire  stopEn125;
  wire  stopEn126;
  wire  stopEn127;
  wire  stopEn128;
  wire  stopEn129;
  wire  stopEn130;
  wire  stopEn131;
  wire  stopEn132;
  wire  stopEn133;
  wire  stopEn134;
  wire  stopEn135;
  wire  stopEn136;
  wire  stopEn137;
  wire  stopEn138;
  wire  stopEn139;
  wire  stopEn140;
  wire  stopEn141;
  wire  stopEn142;
  wire  stopEn143;
  wire  stopEn144;
  wire  stopEn145;
  wire  stopEn146;
  wire  stopEn147;
  wire  stopEn148;
  wire  stopEn149;
  wire  stopEn150;
  wire  stopEn151;
  wire  stopEn152;
  wire  stopEn153;
  wire  stopEn154;
  wire  stopEn155;
  wire  stopEn156;
  wire  stopEn157;
  wire  stopEn158;
  wire  stopEn159;
  wire  stopEn160;
  wire  stopEn161;
  wire  stopEn162;
  wire  stopEn163;
  wire  stopEn164;
  wire  stopEn165;
  wire  stopEn166;
  wire  stopEn167;
  wire  stopEn168;
  wire  stopEn169;
  wire  stopEn170;
  wire  stopEn171;
  wire  stopEn172;
  wire  stopEn173;
  wire  stopEn174;
  wire  stopEn175;
  wire  TLMonitor_66_or63;
  wire  TLMonitor_66_or130;
  wire  TLMonitor_66_or64;
  wire  TLMonitor_66_or31;
  wire  TLMonitor_66_or132;
  wire  TLMonitor_66_or65;
  wire  TLMonitor_66_or134;
  wire  TLMonitor_66_or66;
  wire  TLMonitor_66_or32;
  wire  TLMonitor_66_or15;
  wire  TLMonitor_66_or67;
  wire  TLMonitor_66_or138;
  wire  TLMonitor_66_or68;
  wire  TLMonitor_66_or33;
  wire  TLMonitor_66_or140;
  wire  TLMonitor_66_or69;
  wire  TLMonitor_66_or142;
  wire  TLMonitor_66_or70;
  wire  TLMonitor_66_or34;
  wire  TLMonitor_66_or16;
  wire  TLMonitor_66_or7;
  wire  TLMonitor_66_or71;
  wire  TLMonitor_66_or146;
  wire  TLMonitor_66_or72;
  wire  TLMonitor_66_or35;
  wire  TLMonitor_66_or148;
  wire  TLMonitor_66_or73;
  wire  TLMonitor_66_or150;
  wire  TLMonitor_66_or74;
  wire  TLMonitor_66_or36;
  wire  TLMonitor_66_or17;
  wire  TLMonitor_66_or75;
  wire  TLMonitor_66_or154;
  wire  TLMonitor_66_or76;
  wire  TLMonitor_66_or37;
  wire  TLMonitor_66_or156;
  wire  TLMonitor_66_or77;
  wire  TLMonitor_66_or158;
  wire  TLMonitor_66_or78;
  wire  TLMonitor_66_or38;
  wire  TLMonitor_66_or18;
  wire  TLMonitor_66_or8;
  wire  TLMonitor_66_or3;
  wire  TLMonitor_66_or79;
  wire  TLMonitor_66_or162;
  wire  TLMonitor_66_or80;
  wire  TLMonitor_66_or39;
  wire  TLMonitor_66_or164;
  wire  TLMonitor_66_or81;
  wire  TLMonitor_66_or166;
  wire  TLMonitor_66_or82;
  wire  TLMonitor_66_or40;
  wire  TLMonitor_66_or19;
  wire  TLMonitor_66_or83;
  wire  TLMonitor_66_or170;
  wire  TLMonitor_66_or84;
  wire  TLMonitor_66_or41;
  wire  TLMonitor_66_or172;
  wire  TLMonitor_66_or85;
  wire  TLMonitor_66_or174;
  wire  TLMonitor_66_or86;
  wire  TLMonitor_66_or42;
  wire  TLMonitor_66_or20;
  wire  TLMonitor_66_or9;
  wire  TLMonitor_66_or87;
  wire  TLMonitor_66_or178;
  wire  TLMonitor_66_or88;
  wire  TLMonitor_66_or43;
  wire  TLMonitor_66_or180;
  wire  TLMonitor_66_or89;
  wire  TLMonitor_66_or182;
  wire  TLMonitor_66_or90;
  wire  TLMonitor_66_or44;
  wire  TLMonitor_66_or21;
  wire  TLMonitor_66_or91;
  wire  TLMonitor_66_or186;
  wire  TLMonitor_66_or92;
  wire  TLMonitor_66_or45;
  wire  TLMonitor_66_or188;
  wire  TLMonitor_66_or93;
  wire  TLMonitor_66_or190;
  wire  TLMonitor_66_or94;
  wire  TLMonitor_66_or46;
  wire  TLMonitor_66_or22;
  wire  TLMonitor_66_or10;
  wire  TLMonitor_66_or4;
  wire  TLMonitor_66_or1;
  wire  TLMonitor_66_or95;
  wire  TLMonitor_66_or194;
  wire  TLMonitor_66_or96;
  wire  TLMonitor_66_or47;
  wire  TLMonitor_66_or196;
  wire  TLMonitor_66_or97;
  wire  TLMonitor_66_or198;
  wire  TLMonitor_66_or98;
  wire  TLMonitor_66_or48;
  wire  TLMonitor_66_or23;
  wire  TLMonitor_66_or99;
  wire  TLMonitor_66_or202;
  wire  TLMonitor_66_or100;
  wire  TLMonitor_66_or49;
  wire  TLMonitor_66_or204;
  wire  TLMonitor_66_or101;
  wire  TLMonitor_66_or206;
  wire  TLMonitor_66_or102;
  wire  TLMonitor_66_or50;
  wire  TLMonitor_66_or24;
  wire  TLMonitor_66_or11;
  wire  TLMonitor_66_or103;
  wire  TLMonitor_66_or210;
  wire  TLMonitor_66_or104;
  wire  TLMonitor_66_or51;
  wire  TLMonitor_66_or212;
  wire  TLMonitor_66_or105;
  wire  TLMonitor_66_or214;
  wire  TLMonitor_66_or106;
  wire  TLMonitor_66_or52;
  wire  TLMonitor_66_or25;
  wire  TLMonitor_66_or107;
  wire  TLMonitor_66_or218;
  wire  TLMonitor_66_or108;
  wire  TLMonitor_66_or53;
  wire  TLMonitor_66_or220;
  wire  TLMonitor_66_or109;
  wire  TLMonitor_66_or222;
  wire  TLMonitor_66_or110;
  wire  TLMonitor_66_or54;
  wire  TLMonitor_66_or26;
  wire  TLMonitor_66_or12;
  wire  TLMonitor_66_or5;
  wire  TLMonitor_66_or111;
  wire  TLMonitor_66_or226;
  wire  TLMonitor_66_or112;
  wire  TLMonitor_66_or55;
  wire  TLMonitor_66_or228;
  wire  TLMonitor_66_or113;
  wire  TLMonitor_66_or230;
  wire  TLMonitor_66_or114;
  wire  TLMonitor_66_or56;
  wire  TLMonitor_66_or27;
  wire  TLMonitor_66_or115;
  wire  TLMonitor_66_or234;
  wire  TLMonitor_66_or116;
  wire  TLMonitor_66_or57;
  wire  TLMonitor_66_or236;
  wire  TLMonitor_66_or117;
  wire  TLMonitor_66_or238;
  wire  TLMonitor_66_or118;
  wire  TLMonitor_66_or58;
  wire  TLMonitor_66_or28;
  wire  TLMonitor_66_or13;
  wire  TLMonitor_66_or119;
  wire  TLMonitor_66_or242;
  wire  TLMonitor_66_or120;
  wire  TLMonitor_66_or59;
  wire  TLMonitor_66_or244;
  wire  TLMonitor_66_or121;
  wire  TLMonitor_66_or246;
  wire  TLMonitor_66_or122;
  wire  TLMonitor_66_or60;
  wire  TLMonitor_66_or29;
  wire  TLMonitor_66_or123;
  wire  TLMonitor_66_or250;
  wire  TLMonitor_66_or124;
  wire  TLMonitor_66_or61;
  wire  TLMonitor_66_or252;
  wire  TLMonitor_66_or125;
  wire  TLMonitor_66_or254;
  wire  TLMonitor_66_or126;
  wire  TLMonitor_66_or62;
  wire  TLMonitor_66_or30;
  wire  TLMonitor_66_or14;
  wire  TLMonitor_66_or6;
  wire  TLMonitor_66_or2;
  wire  TLMonitor_66_or0;
  reg  TLMonitor_66_metaAssert;
  reg [31:0] _RAND_30;
  assign _T_20 = io_in_a_bits_source == 2'h0; // @[Parameters.scala 44:9]
  assign _T_21 = io_in_a_bits_source == 2'h1; // @[Parameters.scala 44:9]
  assign _T_22 = io_in_a_bits_source == 2'h2; // @[Parameters.scala 44:9]
  assign _T_32 = _T_20 | _T_21; // @[Parameters.scala 280:46]
  assign _T_33 = _T_32 | _T_22; // @[Parameters.scala 280:46]
  assign _T_35 = 27'hfff << io_in_a_bits_size; // @[package.scala 185:77]
  assign _GEN_33 = {{20'd0}, ~_T_35[11:0]}; // @[Edges.scala 21:16]
  assign _T_38 = io_in_a_bits_address & _GEN_33; // @[Edges.scala 21:16]
  assign _T_39 = _T_38 == 32'h0; // @[Edges.scala 21:24]
  assign _T_42 = 4'h1 << io_in_a_bits_size[1:0]; // @[OneHot.scala 52:12]
  assign _T_44 = _T_42[2:0] | 3'h1; // @[Misc.scala 206:81]
  assign _T_45 = io_in_a_bits_size >= 4'h3; // @[Misc.scala 210:21]
  assign _T_50 = _T_44[2] & ~io_in_a_bits_address[2]; // @[Misc.scala 219:38]
  assign _T_51 = _T_45 | _T_50; // @[Misc.scala 219:29]
  assign _T_53 = _T_44[2] & io_in_a_bits_address[2]; // @[Misc.scala 219:38]
  assign _T_54 = _T_45 | _T_53; // @[Misc.scala 219:29]
  assign _T_58 = ~io_in_a_bits_address[2] & ~io_in_a_bits_address[1]; // @[Misc.scala 218:27]
  assign _T_59 = _T_44[1] & _T_58; // @[Misc.scala 219:38]
  assign _T_60 = _T_51 | _T_59; // @[Misc.scala 219:29]
  assign _T_61 = ~io_in_a_bits_address[2] & io_in_a_bits_address[1]; // @[Misc.scala 218:27]
  assign _T_62 = _T_44[1] & _T_61; // @[Misc.scala 219:38]
  assign _T_63 = _T_51 | _T_62; // @[Misc.scala 219:29]
  assign _T_64 = io_in_a_bits_address[2] & ~io_in_a_bits_address[1]; // @[Misc.scala 218:27]
  assign _T_65 = _T_44[1] & _T_64; // @[Misc.scala 219:38]
  assign _T_66 = _T_54 | _T_65; // @[Misc.scala 219:29]
  assign _T_67 = io_in_a_bits_address[2] & io_in_a_bits_address[1]; // @[Misc.scala 218:27]
  assign _T_68 = _T_44[1] & _T_67; // @[Misc.scala 219:38]
  assign _T_69 = _T_54 | _T_68; // @[Misc.scala 219:29]
  assign _T_73 = _T_58 & ~io_in_a_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_74 = _T_44[0] & _T_73; // @[Misc.scala 219:38]
  assign _T_75 = _T_60 | _T_74; // @[Misc.scala 219:29]
  assign _T_76 = _T_58 & io_in_a_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_77 = _T_44[0] & _T_76; // @[Misc.scala 219:38]
  assign _T_78 = _T_60 | _T_77; // @[Misc.scala 219:29]
  assign _T_79 = _T_61 & ~io_in_a_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_80 = _T_44[0] & _T_79; // @[Misc.scala 219:38]
  assign _T_81 = _T_63 | _T_80; // @[Misc.scala 219:29]
  assign _T_82 = _T_61 & io_in_a_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_83 = _T_44[0] & _T_82; // @[Misc.scala 219:38]
  assign _T_84 = _T_63 | _T_83; // @[Misc.scala 219:29]
  assign _T_85 = _T_64 & ~io_in_a_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_86 = _T_44[0] & _T_85; // @[Misc.scala 219:38]
  assign _T_87 = _T_66 | _T_86; // @[Misc.scala 219:29]
  assign _T_88 = _T_64 & io_in_a_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_89 = _T_44[0] & _T_88; // @[Misc.scala 219:38]
  assign _T_90 = _T_66 | _T_89; // @[Misc.scala 219:29]
  assign _T_91 = _T_67 & ~io_in_a_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_92 = _T_44[0] & _T_91; // @[Misc.scala 219:38]
  assign _T_93 = _T_69 | _T_92; // @[Misc.scala 219:29]
  assign _T_94 = _T_67 & io_in_a_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_95 = _T_44[0] & _T_94; // @[Misc.scala 219:38]
  assign _T_96 = _T_69 | _T_95; // @[Misc.scala 219:29]
  assign _T_103 = {_T_96,_T_93,_T_90,_T_87,_T_84,_T_81,_T_78,_T_75}; // @[Cat.scala 30:58]
  assign _T_107 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 121:49]
  assign _T_133 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 48:25]
  assign _T_135 = io_in_a_bits_size <= 4'h6; // @[Parameters.scala 90:42]
  assign _T_138 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 121:31]
  assign _T_139 = {1'b0,$signed(_T_138)}; // @[Parameters.scala 121:49]
  assign _T_141 = $signed(_T_139) & -33'sh10000000; // @[Parameters.scala 121:52]
  assign _T_142 = $signed(_T_141) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_143 = _T_135 & _T_142; // @[Parameters.scala 168:56]
  assign _T_145 = io_in_a_bits_address ^ 32'h3000; // @[Parameters.scala 121:31]
  assign _T_146 = {1'b0,$signed(_T_145)}; // @[Parameters.scala 121:49]
  assign _T_148 = $signed(_T_146) & -33'sh1000; // @[Parameters.scala 121:52]
  assign _T_149 = $signed(_T_148) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_150 = io_in_a_bits_address ^ 32'hc000000; // @[Parameters.scala 121:31]
  assign _T_151 = {1'b0,$signed(_T_150)}; // @[Parameters.scala 121:49]
  assign _T_153 = $signed(_T_151) & -33'sh4000000; // @[Parameters.scala 121:52]
  assign _T_154 = $signed(_T_153) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_155 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 121:31]
  assign _T_156 = {1'b0,$signed(_T_155)}; // @[Parameters.scala 121:49]
  assign _T_158 = $signed(_T_156) & -33'sh10000; // @[Parameters.scala 121:52]
  assign _T_159 = $signed(_T_158) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_163 = $signed(_T_107) & -33'sh1000; // @[Parameters.scala 121:52]
  assign _T_164 = $signed(_T_163) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_165 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 121:31]
  assign _T_166 = {1'b0,$signed(_T_165)}; // @[Parameters.scala 121:49]
  assign _T_168 = $signed(_T_166) & -33'sh10000; // @[Parameters.scala 121:52]
  assign _T_169 = $signed(_T_168) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_170 = io_in_a_bits_address ^ 32'h60000000; // @[Parameters.scala 121:31]
  assign _T_171 = {1'b0,$signed(_T_170)}; // @[Parameters.scala 121:49]
  assign _T_173 = $signed(_T_171) & -33'sh20000000; // @[Parameters.scala 121:52]
  assign _T_174 = $signed(_T_173) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_175 = _T_149 | _T_154; // @[Parameters.scala 169:42]
  assign _T_176 = _T_175 | _T_159; // @[Parameters.scala 169:42]
  assign _T_177 = _T_176 | _T_164; // @[Parameters.scala 169:42]
  assign _T_184 = _T_143 | reset; // @[Monitor.scala 49:14]
  assign _T_198 = 4'h6 == io_in_a_bits_size; // @[Parameters.scala 89:48]
  assign _T_200 = _T_20 & _T_198; // @[Mux.scala 19:72]
  assign _T_208 = _T_200 | reset; // @[Monitor.scala 50:14]
  assign _T_211 = _T_33 | reset; // @[Monitor.scala 51:14]
  assign _T_215 = _T_45 | reset; // @[Monitor.scala 52:14]
  assign _T_218 = _T_39 | reset; // @[Monitor.scala 53:14]
  assign _T_220 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 109:27]
  assign _T_222 = _T_220 | reset; // @[Monitor.scala 54:14]
  assign _T_225 = ~io_in_a_bits_mask == 8'h0; // @[Monitor.scala 55:28]
  assign _T_227 = _T_225 | reset; // @[Monitor.scala 55:14]
  assign _T_231 = ~io_in_a_bits_corrupt | reset; // @[Monitor.scala 56:14]
  assign _T_233 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 59:25]
  assign _T_324 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 66:28]
  assign _T_326 = _T_324 | reset; // @[Monitor.scala 66:14]
  assign _T_337 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 71:25]
  assign _T_339 = io_in_a_bits_size <= 4'hc; // @[Parameters.scala 90:42]
  assign _T_347 = _T_339 & _T_149; // @[Parameters.scala 168:56]
  assign _T_382 = _T_154 | _T_159; // @[Parameters.scala 169:42]
  assign _T_383 = _T_382 | _T_164; // @[Parameters.scala 169:42]
  assign _T_384 = _T_383 | _T_169; // @[Parameters.scala 169:42]
  assign _T_385 = _T_384 | _T_142; // @[Parameters.scala 169:42]
  assign _T_386 = _T_385 | _T_174; // @[Parameters.scala 169:42]
  assign _T_387 = _T_135 & _T_386; // @[Parameters.scala 168:56]
  assign _T_389 = _T_347 | _T_387; // @[Parameters.scala 170:30]
  assign _T_391 = _T_389 | reset; // @[Monitor.scala 72:14]
  assign _T_399 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 75:28]
  assign _T_401 = _T_399 | reset; // @[Monitor.scala 75:14]
  assign _T_403 = io_in_a_bits_mask == _T_103; // @[Monitor.scala 76:27]
  assign _T_405 = _T_403 | reset; // @[Monitor.scala 76:14]
  assign _T_411 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 80:25]
  assign _T_448 = _T_383 | _T_142; // @[Parameters.scala 169:42]
  assign _T_449 = _T_135 & _T_448; // @[Parameters.scala 168:56]
  assign _T_451 = io_in_a_bits_size <= 4'h8; // @[Parameters.scala 90:42]
  assign _T_459 = _T_451 & _T_174; // @[Parameters.scala 168:56]
  assign _T_468 = _T_347 | _T_449; // @[Parameters.scala 170:30]
  assign _T_469 = _T_468 | _T_459; // @[Parameters.scala 170:30]
  assign _T_472 = _T_469 | reset; // @[Monitor.scala 81:14]
  assign _T_488 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 88:25]
  assign _T_562 = io_in_a_bits_mask & ~_T_103; // @[Monitor.scala 93:28]
  assign _T_563 = _T_562 == 8'h0; // @[Monitor.scala 93:37]
  assign _T_565 = _T_563 | reset; // @[Monitor.scala 93:14]
  assign _T_567 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 96:25]
  assign _T_569 = io_in_a_bits_size <= 4'h3; // @[Parameters.scala 90:42]
  assign _T_595 = _T_569 & _T_177; // @[Parameters.scala 168:56]
  assign _T_618 = _T_595 | reset; // @[Monitor.scala 97:14]
  assign _T_626 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 139:33]
  assign _T_628 = _T_626 | reset; // @[Monitor.scala 100:14]
  assign _T_634 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 104:25]
  assign _T_693 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 146:30]
  assign _T_695 = _T_693 | reset; // @[Monitor.scala 108:14]
  assign _T_701 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 112:25]
  assign _T_752 = _T_347 | reset; // @[Monitor.scala 113:14]
  assign _T_768 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 43:24]
  assign _T_770 = _T_768 | reset; // @[Monitor.scala 268:12]
  assign _T_772 = io_in_d_bits_source == 2'h0; // @[Parameters.scala 44:9]
  assign _T_773 = io_in_d_bits_source == 2'h1; // @[Parameters.scala 44:9]
  assign _T_774 = io_in_d_bits_source == 2'h2; // @[Parameters.scala 44:9]
  assign _T_784 = _T_772 | _T_773; // @[Parameters.scala 280:46]
  assign _T_785 = _T_784 | _T_774; // @[Parameters.scala 280:46]
  assign _T_787 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 275:25]
  assign _T_789 = _T_785 | reset; // @[Monitor.scala 276:14]
  assign _T_791 = io_in_d_bits_size >= 4'h3; // @[Monitor.scala 277:27]
  assign _T_793 = _T_791 | reset; // @[Monitor.scala 277:14]
  assign _T_795 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 278:28]
  assign _T_797 = _T_795 | reset; // @[Monitor.scala 278:14]
  assign _T_801 = ~io_in_d_bits_corrupt | reset; // @[Monitor.scala 279:14]
  assign _T_805 = ~io_in_d_bits_denied | reset; // @[Monitor.scala 280:14]
  assign _T_807 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 283:25]
  assign _T_818 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 103:26]
  assign _T_820 = _T_818 | reset; // @[Monitor.scala 287:14]
  assign _T_822 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 288:28]
  assign _T_824 = _T_822 | reset; // @[Monitor.scala 288:14]
  assign _T_835 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 293:25]
  assign _T_855 = ~io_in_d_bits_denied | io_in_d_bits_corrupt; // @[Monitor.scala 299:30]
  assign _T_857 = _T_855 | reset; // @[Monitor.scala 299:14]
  assign _T_864 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 303:25]
  assign _T_881 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 311:25]
  assign _T_899 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 319:25]
  assign _T_916 = io_in_b_bits_opcode <= 3'h6; // @[Bundles.scala 41:24]
  assign _T_918 = _T_916 | reset; // @[Monitor.scala 122:12]
  assign _T_920 = io_in_b_bits_source == 2'h0; // @[Parameters.scala 44:9]
  assign _T_923 = {1'b0,$signed(io_in_b_bits_address)}; // @[Parameters.scala 121:49]
  assign _T_928 = io_in_b_bits_source == 2'h1; // @[Parameters.scala 44:9]
  assign _T_936 = io_in_b_bits_source == 2'h2; // @[Parameters.scala 44:9]
  assign _T_949 = io_in_b_bits_address ^ 32'h3000; // @[Parameters.scala 121:31]
  assign _T_950 = {1'b0,$signed(_T_949)}; // @[Parameters.scala 121:49]
  assign _T_952 = $signed(_T_950) & -33'sh1000; // @[Parameters.scala 121:52]
  assign _T_953 = $signed(_T_952) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_954 = io_in_b_bits_address ^ 32'hc000000; // @[Parameters.scala 121:31]
  assign _T_955 = {1'b0,$signed(_T_954)}; // @[Parameters.scala 121:49]
  assign _T_957 = $signed(_T_955) & -33'sh4000000; // @[Parameters.scala 121:52]
  assign _T_958 = $signed(_T_957) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_959 = io_in_b_bits_address ^ 32'h2000000; // @[Parameters.scala 121:31]
  assign _T_960 = {1'b0,$signed(_T_959)}; // @[Parameters.scala 121:49]
  assign _T_962 = $signed(_T_960) & -33'sh10000; // @[Parameters.scala 121:52]
  assign _T_963 = $signed(_T_962) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_967 = $signed(_T_923) & -33'sh1000; // @[Parameters.scala 121:52]
  assign _T_968 = $signed(_T_967) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_969 = io_in_b_bits_address ^ 32'h10000; // @[Parameters.scala 121:31]
  assign _T_970 = {1'b0,$signed(_T_969)}; // @[Parameters.scala 121:49]
  assign _T_972 = $signed(_T_970) & -33'sh10000; // @[Parameters.scala 121:52]
  assign _T_973 = $signed(_T_972) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_974 = io_in_b_bits_address ^ 32'h80000000; // @[Parameters.scala 121:31]
  assign _T_975 = {1'b0,$signed(_T_974)}; // @[Parameters.scala 121:49]
  assign _T_977 = $signed(_T_975) & -33'sh10000000; // @[Parameters.scala 121:52]
  assign _T_978 = $signed(_T_977) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_979 = io_in_b_bits_address ^ 32'h60000000; // @[Parameters.scala 121:31]
  assign _T_980 = {1'b0,$signed(_T_979)}; // @[Parameters.scala 121:49]
  assign _T_982 = $signed(_T_980) & -33'sh20000000; // @[Parameters.scala 121:52]
  assign _T_983 = $signed(_T_982) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_997 = _T_953 | _T_958; // @[Parameters.scala 155:64]
  assign _T_998 = _T_997 | _T_963; // @[Parameters.scala 155:64]
  assign _T_999 = _T_998 | _T_968; // @[Parameters.scala 155:64]
  assign _T_1000 = _T_999 | _T_973; // @[Parameters.scala 155:64]
  assign _T_1001 = _T_1000 | _T_978; // @[Parameters.scala 155:64]
  assign _T_1002 = _T_1001 | _T_983; // @[Parameters.scala 155:64]
  assign _T_1004 = 27'hfff << io_in_b_bits_size; // @[package.scala 185:77]
  assign _GEN_34 = {{20'd0}, ~_T_1004[11:0]}; // @[Edges.scala 21:16]
  assign _T_1007 = io_in_b_bits_address & _GEN_34; // @[Edges.scala 21:16]
  assign _T_1008 = _T_1007 == 32'h0; // @[Edges.scala 21:24]
  assign _T_1011 = 4'h1 << io_in_b_bits_size[1:0]; // @[OneHot.scala 52:12]
  assign _T_1013 = _T_1011[2:0] | 3'h1; // @[Misc.scala 206:81]
  assign _T_1014 = io_in_b_bits_size >= 4'h3; // @[Misc.scala 210:21]
  assign _T_1019 = _T_1013[2] & ~io_in_b_bits_address[2]; // @[Misc.scala 219:38]
  assign _T_1020 = _T_1014 | _T_1019; // @[Misc.scala 219:29]
  assign _T_1022 = _T_1013[2] & io_in_b_bits_address[2]; // @[Misc.scala 219:38]
  assign _T_1023 = _T_1014 | _T_1022; // @[Misc.scala 219:29]
  assign _T_1027 = ~io_in_b_bits_address[2] & ~io_in_b_bits_address[1]; // @[Misc.scala 218:27]
  assign _T_1028 = _T_1013[1] & _T_1027; // @[Misc.scala 219:38]
  assign _T_1029 = _T_1020 | _T_1028; // @[Misc.scala 219:29]
  assign _T_1030 = ~io_in_b_bits_address[2] & io_in_b_bits_address[1]; // @[Misc.scala 218:27]
  assign _T_1031 = _T_1013[1] & _T_1030; // @[Misc.scala 219:38]
  assign _T_1032 = _T_1020 | _T_1031; // @[Misc.scala 219:29]
  assign _T_1033 = io_in_b_bits_address[2] & ~io_in_b_bits_address[1]; // @[Misc.scala 218:27]
  assign _T_1034 = _T_1013[1] & _T_1033; // @[Misc.scala 219:38]
  assign _T_1035 = _T_1023 | _T_1034; // @[Misc.scala 219:29]
  assign _T_1036 = io_in_b_bits_address[2] & io_in_b_bits_address[1]; // @[Misc.scala 218:27]
  assign _T_1037 = _T_1013[1] & _T_1036; // @[Misc.scala 219:38]
  assign _T_1038 = _T_1023 | _T_1037; // @[Misc.scala 219:29]
  assign _T_1042 = _T_1027 & ~io_in_b_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_1043 = _T_1013[0] & _T_1042; // @[Misc.scala 219:38]
  assign _T_1044 = _T_1029 | _T_1043; // @[Misc.scala 219:29]
  assign _T_1045 = _T_1027 & io_in_b_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_1046 = _T_1013[0] & _T_1045; // @[Misc.scala 219:38]
  assign _T_1047 = _T_1029 | _T_1046; // @[Misc.scala 219:29]
  assign _T_1048 = _T_1030 & ~io_in_b_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_1049 = _T_1013[0] & _T_1048; // @[Misc.scala 219:38]
  assign _T_1050 = _T_1032 | _T_1049; // @[Misc.scala 219:29]
  assign _T_1051 = _T_1030 & io_in_b_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_1052 = _T_1013[0] & _T_1051; // @[Misc.scala 219:38]
  assign _T_1053 = _T_1032 | _T_1052; // @[Misc.scala 219:29]
  assign _T_1054 = _T_1033 & ~io_in_b_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_1055 = _T_1013[0] & _T_1054; // @[Misc.scala 219:38]
  assign _T_1056 = _T_1035 | _T_1055; // @[Misc.scala 219:29]
  assign _T_1057 = _T_1033 & io_in_b_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_1058 = _T_1013[0] & _T_1057; // @[Misc.scala 219:38]
  assign _T_1059 = _T_1035 | _T_1058; // @[Misc.scala 219:29]
  assign _T_1060 = _T_1036 & ~io_in_b_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_1061 = _T_1013[0] & _T_1060; // @[Misc.scala 219:38]
  assign _T_1062 = _T_1038 | _T_1061; // @[Misc.scala 219:29]
  assign _T_1063 = _T_1036 & io_in_b_bits_address[0]; // @[Misc.scala 218:27]
  assign _T_1064 = _T_1013[0] & _T_1063; // @[Misc.scala 219:38]
  assign _T_1065 = _T_1038 | _T_1064; // @[Misc.scala 219:29]
  assign _T_1072 = {_T_1065,_T_1062,_T_1059,_T_1056,_T_1053,_T_1050,_T_1047,_T_1044}; // @[Cat.scala 30:58]
  assign _T_1088 = _T_936 ? 2'h2 : 2'h0; // @[Mux.scala 19:72]
  assign _GEN_35 = {{1'd0}, _T_928}; // @[Mux.scala 19:72]
  assign _T_1090 = _GEN_35 | _T_1088; // @[Mux.scala 19:72]
  assign _T_1093 = _T_1090 == io_in_b_bits_source; // @[Monitor.scala 130:117]
  assign _T_1094 = io_in_b_bits_opcode == 3'h6; // @[Monitor.scala 132:25]
  assign _T_1107 = 4'h6 == io_in_b_bits_size; // @[Parameters.scala 89:48]
  assign _T_1109 = _T_920 & _T_1107; // @[Mux.scala 19:72]
  assign _T_1117 = _T_1109 | reset; // @[Monitor.scala 133:14]
  assign _T_1120 = _T_1002 | reset; // @[Monitor.scala 134:14]
  assign _T_1123 = _T_1093 | reset; // @[Monitor.scala 135:14]
  assign _T_1126 = _T_1008 | reset; // @[Monitor.scala 136:14]
  assign _T_1128 = io_in_b_bits_param <= 2'h2; // @[Bundles.scala 103:26]
  assign _T_1130 = _T_1128 | reset; // @[Monitor.scala 137:14]
  assign _T_1132 = io_in_b_bits_mask == _T_1072; // @[Monitor.scala 138:27]
  assign _T_1134 = _T_1132 | reset; // @[Monitor.scala 138:14]
  assign _T_1138 = ~io_in_b_bits_corrupt | reset; // @[Monitor.scala 139:14]
  assign _T_1140 = io_in_b_bits_opcode == 3'h4; // @[Monitor.scala 142:25]
  assign _T_1153 = io_in_b_bits_param == 2'h0; // @[Monitor.scala 147:28]
  assign _T_1155 = _T_1153 | reset; // @[Monitor.scala 147:14]
  assign _T_1165 = io_in_b_bits_opcode == 3'h0; // @[Monitor.scala 152:25]
  assign _T_1186 = io_in_b_bits_opcode == 3'h1; // @[Monitor.scala 161:25]
  assign _T_1204 = io_in_b_bits_mask & ~_T_1072; // @[Monitor.scala 167:28]
  assign _T_1205 = _T_1204 == 8'h0; // @[Monitor.scala 167:37]
  assign _T_1207 = _T_1205 | reset; // @[Monitor.scala 167:14]
  assign _T_1209 = io_in_b_bits_opcode == 3'h2; // @[Monitor.scala 170:25]
  assign _T_1230 = io_in_b_bits_opcode == 3'h3; // @[Monitor.scala 179:25]
  assign _T_1251 = io_in_b_bits_opcode == 3'h5; // @[Monitor.scala 188:25]
  assign _T_1276 = io_in_c_bits_source == 2'h0; // @[Parameters.scala 44:9]
  assign _T_1277 = io_in_c_bits_source == 2'h1; // @[Parameters.scala 44:9]
  assign _T_1278 = io_in_c_bits_source == 2'h2; // @[Parameters.scala 44:9]
  assign _T_1288 = _T_1276 | _T_1277; // @[Parameters.scala 280:46]
  assign _T_1289 = _T_1288 | _T_1278; // @[Parameters.scala 280:46]
  assign _T_1291 = 27'hfff << io_in_c_bits_size; // @[package.scala 185:77]
  assign _GEN_36 = {{20'd0}, ~_T_1291[11:0]}; // @[Edges.scala 21:16]
  assign _T_1294 = io_in_c_bits_address & _GEN_36; // @[Edges.scala 21:16]
  assign _T_1295 = _T_1294 == 32'h0; // @[Edges.scala 21:24]
  assign _T_1296 = io_in_c_bits_address ^ 32'h3000; // @[Parameters.scala 121:31]
  assign _T_1297 = {1'b0,$signed(_T_1296)}; // @[Parameters.scala 121:49]
  assign _T_1299 = $signed(_T_1297) & -33'sh1000; // @[Parameters.scala 121:52]
  assign _T_1300 = $signed(_T_1299) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_1301 = io_in_c_bits_address ^ 32'hc000000; // @[Parameters.scala 121:31]
  assign _T_1302 = {1'b0,$signed(_T_1301)}; // @[Parameters.scala 121:49]
  assign _T_1304 = $signed(_T_1302) & -33'sh4000000; // @[Parameters.scala 121:52]
  assign _T_1305 = $signed(_T_1304) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_1306 = io_in_c_bits_address ^ 32'h2000000; // @[Parameters.scala 121:31]
  assign _T_1307 = {1'b0,$signed(_T_1306)}; // @[Parameters.scala 121:49]
  assign _T_1309 = $signed(_T_1307) & -33'sh10000; // @[Parameters.scala 121:52]
  assign _T_1310 = $signed(_T_1309) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_1312 = {1'b0,$signed(io_in_c_bits_address)}; // @[Parameters.scala 121:49]
  assign _T_1314 = $signed(_T_1312) & -33'sh1000; // @[Parameters.scala 121:52]
  assign _T_1315 = $signed(_T_1314) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_1316 = io_in_c_bits_address ^ 32'h10000; // @[Parameters.scala 121:31]
  assign _T_1317 = {1'b0,$signed(_T_1316)}; // @[Parameters.scala 121:49]
  assign _T_1319 = $signed(_T_1317) & -33'sh10000; // @[Parameters.scala 121:52]
  assign _T_1320 = $signed(_T_1319) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_1321 = io_in_c_bits_address ^ 32'h80000000; // @[Parameters.scala 121:31]
  assign _T_1322 = {1'b0,$signed(_T_1321)}; // @[Parameters.scala 121:49]
  assign _T_1324 = $signed(_T_1322) & -33'sh10000000; // @[Parameters.scala 121:52]
  assign _T_1325 = $signed(_T_1324) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_1326 = io_in_c_bits_address ^ 32'h60000000; // @[Parameters.scala 121:31]
  assign _T_1327 = {1'b0,$signed(_T_1326)}; // @[Parameters.scala 121:49]
  assign _T_1329 = $signed(_T_1327) & -33'sh20000000; // @[Parameters.scala 121:52]
  assign _T_1330 = $signed(_T_1329) == 33'sh0; // @[Parameters.scala 121:67]
  assign _T_1344 = _T_1300 | _T_1305; // @[Parameters.scala 155:64]
  assign _T_1345 = _T_1344 | _T_1310; // @[Parameters.scala 155:64]
  assign _T_1346 = _T_1345 | _T_1315; // @[Parameters.scala 155:64]
  assign _T_1347 = _T_1346 | _T_1320; // @[Parameters.scala 155:64]
  assign _T_1348 = _T_1347 | _T_1325; // @[Parameters.scala 155:64]
  assign _T_1349 = _T_1348 | _T_1330; // @[Parameters.scala 155:64]
  assign _T_1379 = io_in_c_bits_opcode == 3'h4; // @[Monitor.scala 207:25]
  assign _T_1381 = _T_1349 | reset; // @[Monitor.scala 208:14]
  assign _T_1384 = _T_1289 | reset; // @[Monitor.scala 209:14]
  assign _T_1386 = io_in_c_bits_size >= 4'h3; // @[Monitor.scala 210:27]
  assign _T_1388 = _T_1386 | reset; // @[Monitor.scala 210:14]
  assign _T_1391 = _T_1295 | reset; // @[Monitor.scala 211:14]
  assign _T_1393 = io_in_c_bits_param <= 3'h5; // @[Bundles.scala 121:29]
  assign _T_1395 = _T_1393 | reset; // @[Monitor.scala 212:14]
  assign _T_1401 = io_in_c_bits_opcode == 3'h5; // @[Monitor.scala 216:25]
  assign _T_1419 = io_in_c_bits_opcode == 3'h6; // @[Monitor.scala 224:25]
  assign _T_1421 = io_in_c_bits_size <= 4'h6; // @[Parameters.scala 90:42]
  assign _T_1429 = _T_1421 & _T_1325; // @[Parameters.scala 168:56]
  assign _T_1470 = _T_1429 | reset; // @[Monitor.scala 225:14]
  assign _T_1484 = 4'h6 == io_in_c_bits_size; // @[Parameters.scala 89:48]
  assign _T_1486 = _T_1276 & _T_1484; // @[Mux.scala 19:72]
  assign _T_1494 = _T_1486 | reset; // @[Monitor.scala 226:14]
  assign _T_1506 = io_in_c_bits_param <= 3'h2; // @[Bundles.scala 115:29]
  assign _T_1508 = _T_1506 | reset; // @[Monitor.scala 230:14]
  assign _T_1514 = io_in_c_bits_opcode == 3'h7; // @[Monitor.scala 234:25]
  assign _T_1605 = io_in_c_bits_opcode == 3'h0; // @[Monitor.scala 243:25]
  assign _T_1615 = io_in_c_bits_param == 3'h0; // @[Monitor.scala 247:28]
  assign _T_1617 = _T_1615 | reset; // @[Monitor.scala 247:14]
  assign _T_1623 = io_in_c_bits_opcode == 3'h1; // @[Monitor.scala 251:25]
  assign _T_1637 = io_in_c_bits_opcode == 3'h2; // @[Monitor.scala 258:25]
  assign _T_1659 = io_in_a_ready & io_in_a_valid; // @[Bundles.scala 277:22]
  assign _T_1664 = ~_T_35[11:3]; // @[Edges.scala 220:59]
  assign _T_1672 = _T_1669 - 9'h1; // @[Edges.scala 230:28]
  assign _T_1673 = _T_1669 == 9'h0; // @[Edges.scala 231:25]
  assign _T_1692 = io_in_a_valid & ~_T_1673; // @[Monitor.scala 354:19]
  assign _T_1693 = io_in_a_bits_opcode == _T_1682; // @[Monitor.scala 355:29]
  assign _T_1695 = _T_1693 | reset; // @[Monitor.scala 355:14]
  assign _T_1697 = io_in_a_bits_param == _T_1684; // @[Monitor.scala 356:29]
  assign _T_1699 = _T_1697 | reset; // @[Monitor.scala 356:14]
  assign _T_1701 = io_in_a_bits_size == _T_1686; // @[Monitor.scala 357:29]
  assign _T_1703 = _T_1701 | reset; // @[Monitor.scala 357:14]
  assign _T_1705 = io_in_a_bits_source == _T_1688; // @[Monitor.scala 358:29]
  assign _T_1707 = _T_1705 | reset; // @[Monitor.scala 358:14]
  assign _T_1709 = io_in_a_bits_address == _T_1690; // @[Monitor.scala 359:29]
  assign _T_1711 = _T_1709 | reset; // @[Monitor.scala 359:14]
  assign _T_1714 = _T_1659 & _T_1673; // @[Monitor.scala 361:20]
  assign _T_1715 = io_in_d_ready & io_in_d_valid; // @[Bundles.scala 277:22]
  assign _T_1717 = 27'hfff << io_in_d_bits_size; // @[package.scala 185:77]
  assign _T_1720 = ~_T_1717[11:3]; // @[Edges.scala 220:59]
  assign _T_1727 = _T_1724 - 9'h1; // @[Edges.scala 230:28]
  assign _T_1728 = _T_1724 == 9'h0; // @[Edges.scala 231:25]
  assign _T_1749 = io_in_d_valid & ~_T_1728; // @[Monitor.scala 424:19]
  assign _T_1750 = io_in_d_bits_opcode == _T_1737; // @[Monitor.scala 425:29]
  assign _T_1752 = _T_1750 | reset; // @[Monitor.scala 425:14]
  assign _T_1754 = io_in_d_bits_param == _T_1739; // @[Monitor.scala 426:29]
  assign _T_1756 = _T_1754 | reset; // @[Monitor.scala 426:14]
  assign _T_1758 = io_in_d_bits_size == _T_1741; // @[Monitor.scala 427:29]
  assign _T_1760 = _T_1758 | reset; // @[Monitor.scala 427:14]
  assign _T_1762 = io_in_d_bits_source == _T_1743; // @[Monitor.scala 428:29]
  assign _T_1764 = _T_1762 | reset; // @[Monitor.scala 428:14]
  assign _T_1766 = io_in_d_bits_sink == _T_1745; // @[Monitor.scala 429:29]
  assign _T_1768 = _T_1766 | reset; // @[Monitor.scala 429:14]
  assign _T_1770 = io_in_d_bits_denied == _T_1747; // @[Monitor.scala 430:29]
  assign _T_1772 = _T_1770 | reset; // @[Monitor.scala 430:14]
  assign _T_1775 = _T_1715 & _T_1728; // @[Monitor.scala 432:20]
  assign _T_1776 = io_in_b_ready & io_in_b_valid; // @[Bundles.scala 277:22]
  assign _T_1789 = _T_1786 - 9'h1; // @[Edges.scala 230:28]
  assign _T_1790 = _T_1786 == 9'h0; // @[Edges.scala 231:25]
  assign _T_1809 = io_in_b_valid & ~_T_1790; // @[Monitor.scala 377:19]
  assign _T_1810 = io_in_b_bits_opcode == _T_1799; // @[Monitor.scala 378:29]
  assign _T_1812 = _T_1810 | reset; // @[Monitor.scala 378:14]
  assign _T_1814 = io_in_b_bits_param == _T_1801; // @[Monitor.scala 379:29]
  assign _T_1816 = _T_1814 | reset; // @[Monitor.scala 379:14]
  assign _T_1818 = io_in_b_bits_size == _T_1803; // @[Monitor.scala 380:29]
  assign _T_1820 = _T_1818 | reset; // @[Monitor.scala 380:14]
  assign _T_1822 = io_in_b_bits_source == _T_1805; // @[Monitor.scala 381:29]
  assign _T_1824 = _T_1822 | reset; // @[Monitor.scala 381:14]
  assign _T_1826 = io_in_b_bits_address == _T_1807; // @[Monitor.scala 382:29]
  assign _T_1828 = _T_1826 | reset; // @[Monitor.scala 382:14]
  assign _T_1831 = _T_1776 & _T_1790; // @[Monitor.scala 384:20]
  assign _T_1832 = io_in_c_ready & io_in_c_valid; // @[Bundles.scala 277:22]
  assign _T_1837 = ~_T_1291[11:3]; // @[Edges.scala 220:59]
  assign _T_1844 = _T_1841 - 9'h1; // @[Edges.scala 230:28]
  assign _T_1845 = _T_1841 == 9'h0; // @[Edges.scala 231:25]
  assign _T_1864 = io_in_c_valid & ~_T_1845; // @[Monitor.scala 400:19]
  assign _T_1865 = io_in_c_bits_opcode == _T_1854; // @[Monitor.scala 401:29]
  assign _T_1867 = _T_1865 | reset; // @[Monitor.scala 401:14]
  assign _T_1869 = io_in_c_bits_param == _T_1856; // @[Monitor.scala 402:29]
  assign _T_1871 = _T_1869 | reset; // @[Monitor.scala 402:14]
  assign _T_1873 = io_in_c_bits_size == _T_1858; // @[Monitor.scala 403:29]
  assign _T_1875 = _T_1873 | reset; // @[Monitor.scala 403:14]
  assign _T_1877 = io_in_c_bits_source == _T_1860; // @[Monitor.scala 404:29]
  assign _T_1879 = _T_1877 | reset; // @[Monitor.scala 404:14]
  assign _T_1881 = io_in_c_bits_address == _T_1862; // @[Monitor.scala 405:29]
  assign _T_1883 = _T_1881 | reset; // @[Monitor.scala 405:14]
  assign _T_1886 = _T_1832 & _T_1845; // @[Monitor.scala 407:20]
  assign _T_1902 = _T_1899 - 9'h1; // @[Edges.scala 230:28]
  assign _T_1903 = _T_1899 == 9'h0; // @[Edges.scala 231:25]
  assign _T_1923 = _T_1920 - 9'h1; // @[Edges.scala 230:28]
  assign _T_1924 = _T_1920 == 9'h0; // @[Edges.scala 231:25]
  assign _T_1935 = _T_1659 & _T_1903; // @[Monitor.scala 458:27]
  assign _T_1937 = 4'h1 << io_in_a_bits_source; // @[OneHot.scala 45:35]
  assign _T_1938 = _T_1888 >> io_in_a_bits_source; // @[Monitor.scala 460:23]
  assign _T_1942 = ~_T_1938[0] | reset; // @[Monitor.scala 460:13]
  assign _GEN_27 = _T_1935 ? _T_1937 : 4'h0; // @[Monitor.scala 458:72]
  assign _T_1948 = _T_1715 & _T_1924; // @[Monitor.scala 465:27]
  assign _T_1951 = _T_1948 & ~_T_787; // @[Monitor.scala 465:72]
  assign _T_1952 = 4'h1 << io_in_d_bits_source; // @[OneHot.scala 45:35]
  assign _T_1953 = _GEN_27[2:0] | _T_1888; // @[Monitor.scala 467:21]
  assign _T_1954 = _T_1953 >> io_in_d_bits_source; // @[Monitor.scala 467:32]
  assign _T_1957 = _T_1954[0] | reset; // @[Monitor.scala 467:13]
  assign _GEN_28 = _T_1951 ? _T_1952 : 4'h0; // @[Monitor.scala 465:91]
  assign _T_1959 = _GEN_27[2:0] != _GEN_28[2:0]; // @[Monitor.scala 471:20]
  assign _T_1960 = _GEN_27[2:0] != 3'h0; // @[Monitor.scala 471:40]
  assign _T_1962 = _T_1959 | ~_T_1960; // @[Monitor.scala 471:30]
  assign _T_1964 = _T_1962 | reset; // @[Monitor.scala 471:13]
  assign _T_1966 = _T_1888 | _GEN_27[2:0]; // @[Monitor.scala 474:27]
  assign _T_1968 = _T_1966 & ~_GEN_28[2:0]; // @[Monitor.scala 474:36]
  assign _T_1999 = _T_1996 - 9'h1; // @[Edges.scala 230:28]
  assign _T_2000 = _T_1996 == 9'h0; // @[Edges.scala 231:25]
  assign _T_2011 = _T_1715 & _T_2000; // @[Monitor.scala 492:27]
  assign _T_2015 = io_in_d_bits_opcode[2] & ~io_in_d_bits_opcode[1]; // @[Edges.scala 71:40]
  assign _T_2016 = _T_2011 & _T_2015; // @[Monitor.scala 492:38]
  assign _T_2017 = 4'h1 << io_in_d_bits_sink; // @[OneHot.scala 45:35]
  assign _T_2018 = _T_1986 >> io_in_d_bits_sink; // @[Monitor.scala 494:23]
  assign _T_2022 = ~_T_2018[0] | reset; // @[Monitor.scala 494:13]
  assign _GEN_31 = _T_2016 ? _T_2017 : 4'h0; // @[Monitor.scala 492:72]
  assign _T_2026 = io_in_e_ready & io_in_e_valid; // @[Bundles.scala 277:22]
  assign _T_2029 = 4'h1 << io_in_e_bits_sink; // @[OneHot.scala 45:35]
  assign _T_2030 = _GEN_31 | _T_1986; // @[Monitor.scala 500:21]
  assign _T_2031 = _T_2030 >> io_in_e_bits_sink; // @[Monitor.scala 500:32]
  assign _T_2034 = _T_2031[0] | reset; // @[Monitor.scala 500:13]
  assign _GEN_32 = _T_2026 ? _T_2029 : 4'h0; // @[Monitor.scala 498:73]
  assign _T_2036 = _T_1986 | _GEN_31; // @[Monitor.scala 505:27]
  assign _T_2038 = _T_2036 & ~_GEN_32; // @[Monitor.scala 505:36]
  assign _GEN_37 = io_in_a_valid & _T_133; // @[Monitor.scala 49:14]
  assign _GEN_53 = io_in_a_valid & _T_233; // @[Monitor.scala 60:14]
  assign _GEN_71 = io_in_a_valid & _T_337; // @[Monitor.scala 72:14]
  assign _GEN_83 = io_in_a_valid & _T_411; // @[Monitor.scala 81:14]
  assign _GEN_93 = io_in_a_valid & _T_488; // @[Monitor.scala 89:14]
  assign _GEN_103 = io_in_a_valid & _T_567; // @[Monitor.scala 97:14]
  assign _GEN_113 = io_in_a_valid & _T_634; // @[Monitor.scala 105:14]
  assign _GEN_123 = io_in_a_valid & _T_701; // @[Monitor.scala 113:14]
  assign _GEN_133 = io_in_d_valid & _T_787; // @[Monitor.scala 276:14]
  assign _GEN_143 = io_in_d_valid & _T_807; // @[Monitor.scala 284:14]
  assign _GEN_153 = io_in_d_valid & _T_835; // @[Monitor.scala 294:14]
  assign _GEN_163 = io_in_d_valid & _T_864; // @[Monitor.scala 304:14]
  assign _GEN_169 = io_in_d_valid & _T_881; // @[Monitor.scala 312:14]
  assign _GEN_175 = io_in_d_valid & _T_899; // @[Monitor.scala 320:14]
  assign _GEN_181 = io_in_b_valid & _T_1094; // @[Monitor.scala 133:14]
  assign _GEN_195 = io_in_b_valid & _T_1140; // @[Monitor.scala 143:14]
  assign _GEN_209 = io_in_b_valid & _T_1165; // @[Monitor.scala 153:14]
  assign _GEN_221 = io_in_b_valid & _T_1186; // @[Monitor.scala 162:14]
  assign _GEN_233 = io_in_b_valid & _T_1209; // @[Monitor.scala 171:14]
  assign _GEN_243 = io_in_b_valid & _T_1230; // @[Monitor.scala 180:14]
  assign _GEN_253 = io_in_b_valid & _T_1251; // @[Monitor.scala 189:14]
  assign _GEN_265 = io_in_c_valid & _T_1379; // @[Monitor.scala 208:14]
  assign _GEN_275 = io_in_c_valid & _T_1401; // @[Monitor.scala 217:14]
  assign _GEN_285 = io_in_c_valid & _T_1419; // @[Monitor.scala 225:14]
  assign _GEN_297 = io_in_c_valid & _T_1514; // @[Monitor.scala 235:14]
  assign _GEN_309 = io_in_c_valid & _T_1605; // @[Monitor.scala 244:14]
  assign _GEN_317 = io_in_c_valid & _T_1623; // @[Monitor.scala 252:14]
  assign _GEN_325 = io_in_c_valid & _T_1637; // @[Monitor.scala 259:14]
  assign TLMonitor_66_covSum = 30'h0;
  assign io_covSum = TLMonitor_66_covSum;
  assign stopEn0 = _GEN_37 & ~_T_184;
  assign stopEn1 = _GEN_37 & ~_T_208;
  assign stopEn2 = _GEN_37 & ~_T_211;
  assign stopEn3 = _GEN_37 & ~_T_215;
  assign stopEn4 = _GEN_37 & ~_T_218;
  assign stopEn5 = _GEN_37 & ~_T_222;
  assign stopEn6 = _GEN_37 & ~_T_227;
  assign stopEn7 = _GEN_37 & ~_T_231;
  assign stopEn8 = _GEN_53 & ~_T_184;
  assign stopEn9 = _GEN_53 & ~_T_208;
  assign stopEn10 = _GEN_53 & ~_T_211;
  assign stopEn11 = _GEN_53 & ~_T_215;
  assign stopEn12 = _GEN_53 & ~_T_218;
  assign stopEn13 = _GEN_53 & ~_T_222;
  assign stopEn14 = _GEN_53 & ~_T_326;
  assign stopEn15 = _GEN_53 & ~_T_227;
  assign stopEn16 = _GEN_53 & ~_T_231;
  assign stopEn17 = _GEN_71 & ~_T_391;
  assign stopEn18 = _GEN_71 & ~_T_211;
  assign stopEn19 = _GEN_71 & ~_T_218;
  assign stopEn20 = _GEN_71 & ~_T_401;
  assign stopEn21 = _GEN_71 & ~_T_405;
  assign stopEn22 = _GEN_71 & ~_T_231;
  assign stopEn23 = _GEN_83 & ~_T_472;
  assign stopEn24 = _GEN_83 & ~_T_211;
  assign stopEn25 = _GEN_83 & ~_T_218;
  assign stopEn26 = _GEN_83 & ~_T_401;
  assign stopEn27 = _GEN_83 & ~_T_405;
  assign stopEn28 = _GEN_93 & ~_T_472;
  assign stopEn29 = _GEN_93 & ~_T_211;
  assign stopEn30 = _GEN_93 & ~_T_218;
  assign stopEn31 = _GEN_93 & ~_T_401;
  assign stopEn32 = _GEN_93 & ~_T_565;
  assign stopEn33 = _GEN_103 & ~_T_618;
  assign stopEn34 = _GEN_103 & ~_T_211;
  assign stopEn35 = _GEN_103 & ~_T_218;
  assign stopEn36 = _GEN_103 & ~_T_628;
  assign stopEn37 = _GEN_103 & ~_T_405;
  assign stopEn38 = _GEN_113 & ~_T_618;
  assign stopEn39 = _GEN_113 & ~_T_211;
  assign stopEn40 = _GEN_113 & ~_T_218;
  assign stopEn41 = _GEN_113 & ~_T_695;
  assign stopEn42 = _GEN_113 & ~_T_405;
  assign stopEn43 = _GEN_123 & ~_T_752;
  assign stopEn44 = _GEN_123 & ~_T_211;
  assign stopEn45 = _GEN_123 & ~_T_218;
  assign stopEn46 = _GEN_123 & ~_T_405;
  assign stopEn47 = _GEN_123 & ~_T_231;
  assign stopEn48 = io_in_d_valid & ~_T_770;
  assign stopEn49 = _GEN_133 & ~_T_789;
  assign stopEn50 = _GEN_133 & ~_T_793;
  assign stopEn51 = _GEN_133 & ~_T_797;
  assign stopEn52 = _GEN_133 & ~_T_801;
  assign stopEn53 = _GEN_133 & ~_T_805;
  assign stopEn54 = _GEN_143 & ~_T_789;
  assign stopEn55 = _GEN_143 & ~_T_793;
  assign stopEn56 = _GEN_143 & ~_T_820;
  assign stopEn57 = _GEN_143 & ~_T_824;
  assign stopEn58 = _GEN_143 & ~_T_801;
  assign stopEn59 = _GEN_153 & ~_T_789;
  assign stopEn60 = _GEN_153 & ~_T_793;
  assign stopEn61 = _GEN_153 & ~_T_820;
  assign stopEn62 = _GEN_153 & ~_T_824;
  assign stopEn63 = _GEN_153 & ~_T_857;
  assign stopEn64 = _GEN_163 & ~_T_789;
  assign stopEn65 = _GEN_163 & ~_T_797;
  assign stopEn66 = _GEN_163 & ~_T_801;
  assign stopEn67 = _GEN_169 & ~_T_789;
  assign stopEn68 = _GEN_169 & ~_T_797;
  assign stopEn69 = _GEN_169 & ~_T_857;
  assign stopEn70 = _GEN_175 & ~_T_789;
  assign stopEn71 = _GEN_175 & ~_T_797;
  assign stopEn72 = _GEN_175 & ~_T_801;
  assign stopEn73 = io_in_b_valid & ~_T_918;
  assign stopEn74 = _GEN_181 & ~_T_1117;
  assign stopEn75 = _GEN_181 & ~_T_1120;
  assign stopEn76 = _GEN_181 & ~_T_1123;
  assign stopEn77 = _GEN_181 & ~_T_1126;
  assign stopEn78 = _GEN_181 & ~_T_1130;
  assign stopEn79 = _GEN_181 & ~_T_1134;
  assign stopEn80 = _GEN_181 & ~_T_1138;
  assign stopEn81 = _GEN_195 & ~reset;
  assign stopEn82 = _GEN_195 & ~_T_1120;
  assign stopEn83 = _GEN_195 & ~_T_1123;
  assign stopEn84 = _GEN_195 & ~_T_1126;
  assign stopEn85 = _GEN_195 & ~_T_1155;
  assign stopEn86 = _GEN_195 & ~_T_1134;
  assign stopEn87 = _GEN_195 & ~_T_1138;
  assign stopEn88 = _GEN_209 & ~reset;
  assign stopEn89 = _GEN_209 & ~_T_1120;
  assign stopEn90 = _GEN_209 & ~_T_1123;
  assign stopEn91 = _GEN_209 & ~_T_1126;
  assign stopEn92 = _GEN_209 & ~_T_1155;
  assign stopEn93 = _GEN_209 & ~_T_1134;
  assign stopEn94 = _GEN_221 & ~reset;
  assign stopEn95 = _GEN_221 & ~_T_1120;
  assign stopEn96 = _GEN_221 & ~_T_1123;
  assign stopEn97 = _GEN_221 & ~_T_1126;
  assign stopEn98 = _GEN_221 & ~_T_1155;
  assign stopEn99 = _GEN_221 & ~_T_1207;
  assign stopEn100 = _GEN_233 & ~reset;
  assign stopEn101 = _GEN_233 & ~_T_1120;
  assign stopEn102 = _GEN_233 & ~_T_1123;
  assign stopEn103 = _GEN_233 & ~_T_1126;
  assign stopEn104 = _GEN_233 & ~_T_1134;
  assign stopEn105 = _GEN_243 & ~reset;
  assign stopEn106 = _GEN_243 & ~_T_1120;
  assign stopEn107 = _GEN_243 & ~_T_1123;
  assign stopEn108 = _GEN_243 & ~_T_1126;
  assign stopEn109 = _GEN_243 & ~_T_1134;
  assign stopEn110 = _GEN_253 & ~reset;
  assign stopEn111 = _GEN_253 & ~_T_1120;
  assign stopEn112 = _GEN_253 & ~_T_1123;
  assign stopEn113 = _GEN_253 & ~_T_1126;
  assign stopEn114 = _GEN_253 & ~_T_1134;
  assign stopEn115 = _GEN_253 & ~_T_1138;
  assign stopEn116 = _GEN_265 & ~_T_1381;
  assign stopEn117 = _GEN_265 & ~_T_1384;
  assign stopEn118 = _GEN_265 & ~_T_1388;
  assign stopEn119 = _GEN_265 & ~_T_1391;
  assign stopEn120 = _GEN_265 & ~_T_1395;
  assign stopEn121 = _GEN_275 & ~_T_1381;
  assign stopEn122 = _GEN_275 & ~_T_1384;
  assign stopEn123 = _GEN_275 & ~_T_1388;
  assign stopEn124 = _GEN_275 & ~_T_1391;
  assign stopEn125 = _GEN_275 & ~_T_1395;
  assign stopEn126 = _GEN_285 & ~_T_1470;
  assign stopEn127 = _GEN_285 & ~_T_1494;
  assign stopEn128 = _GEN_285 & ~_T_1384;
  assign stopEn129 = _GEN_285 & ~_T_1388;
  assign stopEn130 = _GEN_285 & ~_T_1391;
  assign stopEn131 = _GEN_285 & ~_T_1508;
  assign stopEn132 = _GEN_297 & ~_T_1470;
  assign stopEn133 = _GEN_297 & ~_T_1494;
  assign stopEn134 = _GEN_297 & ~_T_1384;
  assign stopEn135 = _GEN_297 & ~_T_1388;
  assign stopEn136 = _GEN_297 & ~_T_1391;
  assign stopEn137 = _GEN_297 & ~_T_1508;
  assign stopEn138 = _GEN_309 & ~_T_1381;
  assign stopEn139 = _GEN_309 & ~_T_1384;
  assign stopEn140 = _GEN_309 & ~_T_1391;
  assign stopEn141 = _GEN_309 & ~_T_1617;
  assign stopEn142 = _GEN_317 & ~_T_1381;
  assign stopEn143 = _GEN_317 & ~_T_1384;
  assign stopEn144 = _GEN_317 & ~_T_1391;
  assign stopEn145 = _GEN_317 & ~_T_1617;
  assign stopEn146 = _GEN_325 & ~_T_1381;
  assign stopEn147 = _GEN_325 & ~_T_1384;
  assign stopEn148 = _GEN_325 & ~_T_1391;
  assign stopEn149 = _GEN_325 & ~_T_1617;
  assign stopEn150 = _T_1692 & ~_T_1695;
  assign stopEn151 = _T_1692 & ~_T_1699;
  assign stopEn152 = _T_1692 & ~_T_1703;
  assign stopEn153 = _T_1692 & ~_T_1707;
  assign stopEn154 = _T_1692 & ~_T_1711;
  assign stopEn155 = _T_1749 & ~_T_1752;
  assign stopEn156 = _T_1749 & ~_T_1756;
  assign stopEn157 = _T_1749 & ~_T_1760;
  assign stopEn158 = _T_1749 & ~_T_1764;
  assign stopEn159 = _T_1749 & ~_T_1768;
  assign stopEn160 = _T_1749 & ~_T_1772;
  assign stopEn161 = _T_1809 & ~_T_1812;
  assign stopEn162 = _T_1809 & ~_T_1816;
  assign stopEn163 = _T_1809 & ~_T_1820;
  assign stopEn164 = _T_1809 & ~_T_1824;
  assign stopEn165 = _T_1809 & ~_T_1828;
  assign stopEn166 = _T_1864 & ~_T_1867;
  assign stopEn167 = _T_1864 & ~_T_1871;
  assign stopEn168 = _T_1864 & ~_T_1875;
  assign stopEn169 = _T_1864 & ~_T_1879;
  assign stopEn170 = _T_1864 & ~_T_1883;
  assign stopEn171 = _T_1935 & ~_T_1942;
  assign stopEn172 = _T_1951 & ~_T_1957;
  assign stopEn173 = ~_T_1964;
  assign stopEn174 = _T_2016 & ~_T_2022;
  assign stopEn175 = _T_2026 & ~_T_2034;
  assign TLMonitor_66_or63 = stopEn0 | stopEn1;
  assign TLMonitor_66_or130 = stopEn3 | stopEn4;
  assign TLMonitor_66_or64 = stopEn2 | TLMonitor_66_or130;
  assign TLMonitor_66_or31 = TLMonitor_66_or63 | TLMonitor_66_or64;
  assign TLMonitor_66_or132 = stopEn6 | stopEn7;
  assign TLMonitor_66_or65 = stopEn5 | TLMonitor_66_or132;
  assign TLMonitor_66_or134 = stopEn9 | stopEn10;
  assign TLMonitor_66_or66 = stopEn8 | TLMonitor_66_or134;
  assign TLMonitor_66_or32 = TLMonitor_66_or65 | TLMonitor_66_or66;
  assign TLMonitor_66_or15 = TLMonitor_66_or31 | TLMonitor_66_or32;
  assign TLMonitor_66_or67 = stopEn11 | stopEn12;
  assign TLMonitor_66_or138 = stopEn14 | stopEn15;
  assign TLMonitor_66_or68 = stopEn13 | TLMonitor_66_or138;
  assign TLMonitor_66_or33 = TLMonitor_66_or67 | TLMonitor_66_or68;
  assign TLMonitor_66_or140 = stopEn17 | stopEn18;
  assign TLMonitor_66_or69 = stopEn16 | TLMonitor_66_or140;
  assign TLMonitor_66_or142 = stopEn20 | stopEn21;
  assign TLMonitor_66_or70 = stopEn19 | TLMonitor_66_or142;
  assign TLMonitor_66_or34 = TLMonitor_66_or69 | TLMonitor_66_or70;
  assign TLMonitor_66_or16 = TLMonitor_66_or33 | TLMonitor_66_or34;
  assign TLMonitor_66_or7 = TLMonitor_66_or15 | TLMonitor_66_or16;
  assign TLMonitor_66_or71 = stopEn22 | stopEn23;
  assign TLMonitor_66_or146 = stopEn25 | stopEn26;
  assign TLMonitor_66_or72 = stopEn24 | TLMonitor_66_or146;
  assign TLMonitor_66_or35 = TLMonitor_66_or71 | TLMonitor_66_or72;
  assign TLMonitor_66_or148 = stopEn28 | stopEn29;
  assign TLMonitor_66_or73 = stopEn27 | TLMonitor_66_or148;
  assign TLMonitor_66_or150 = stopEn31 | stopEn32;
  assign TLMonitor_66_or74 = stopEn30 | TLMonitor_66_or150;
  assign TLMonitor_66_or36 = TLMonitor_66_or73 | TLMonitor_66_or74;
  assign TLMonitor_66_or17 = TLMonitor_66_or35 | TLMonitor_66_or36;
  assign TLMonitor_66_or75 = stopEn33 | stopEn34;
  assign TLMonitor_66_or154 = stopEn36 | stopEn37;
  assign TLMonitor_66_or76 = stopEn35 | TLMonitor_66_or154;
  assign TLMonitor_66_or37 = TLMonitor_66_or75 | TLMonitor_66_or76;
  assign TLMonitor_66_or156 = stopEn39 | stopEn40;
  assign TLMonitor_66_or77 = stopEn38 | TLMonitor_66_or156;
  assign TLMonitor_66_or158 = stopEn42 | stopEn43;
  assign TLMonitor_66_or78 = stopEn41 | TLMonitor_66_or158;
  assign TLMonitor_66_or38 = TLMonitor_66_or77 | TLMonitor_66_or78;
  assign TLMonitor_66_or18 = TLMonitor_66_or37 | TLMonitor_66_or38;
  assign TLMonitor_66_or8 = TLMonitor_66_or17 | TLMonitor_66_or18;
  assign TLMonitor_66_or3 = TLMonitor_66_or7 | TLMonitor_66_or8;
  assign TLMonitor_66_or79 = stopEn44 | stopEn45;
  assign TLMonitor_66_or162 = stopEn47 | stopEn48;
  assign TLMonitor_66_or80 = stopEn46 | TLMonitor_66_or162;
  assign TLMonitor_66_or39 = TLMonitor_66_or79 | TLMonitor_66_or80;
  assign TLMonitor_66_or164 = stopEn50 | stopEn51;
  assign TLMonitor_66_or81 = stopEn49 | TLMonitor_66_or164;
  assign TLMonitor_66_or166 = stopEn53 | stopEn54;
  assign TLMonitor_66_or82 = stopEn52 | TLMonitor_66_or166;
  assign TLMonitor_66_or40 = TLMonitor_66_or81 | TLMonitor_66_or82;
  assign TLMonitor_66_or19 = TLMonitor_66_or39 | TLMonitor_66_or40;
  assign TLMonitor_66_or83 = stopEn55 | stopEn56;
  assign TLMonitor_66_or170 = stopEn58 | stopEn59;
  assign TLMonitor_66_or84 = stopEn57 | TLMonitor_66_or170;
  assign TLMonitor_66_or41 = TLMonitor_66_or83 | TLMonitor_66_or84;
  assign TLMonitor_66_or172 = stopEn61 | stopEn62;
  assign TLMonitor_66_or85 = stopEn60 | TLMonitor_66_or172;
  assign TLMonitor_66_or174 = stopEn64 | stopEn65;
  assign TLMonitor_66_or86 = stopEn63 | TLMonitor_66_or174;
  assign TLMonitor_66_or42 = TLMonitor_66_or85 | TLMonitor_66_or86;
  assign TLMonitor_66_or20 = TLMonitor_66_or41 | TLMonitor_66_or42;
  assign TLMonitor_66_or9 = TLMonitor_66_or19 | TLMonitor_66_or20;
  assign TLMonitor_66_or87 = stopEn66 | stopEn67;
  assign TLMonitor_66_or178 = stopEn69 | stopEn70;
  assign TLMonitor_66_or88 = stopEn68 | TLMonitor_66_or178;
  assign TLMonitor_66_or43 = TLMonitor_66_or87 | TLMonitor_66_or88;
  assign TLMonitor_66_or180 = stopEn72 | stopEn73;
  assign TLMonitor_66_or89 = stopEn71 | TLMonitor_66_or180;
  assign TLMonitor_66_or182 = stopEn75 | stopEn76;
  assign TLMonitor_66_or90 = stopEn74 | TLMonitor_66_or182;
  assign TLMonitor_66_or44 = TLMonitor_66_or89 | TLMonitor_66_or90;
  assign TLMonitor_66_or21 = TLMonitor_66_or43 | TLMonitor_66_or44;
  assign TLMonitor_66_or91 = stopEn77 | stopEn78;
  assign TLMonitor_66_or186 = stopEn80 | stopEn81;
  assign TLMonitor_66_or92 = stopEn79 | TLMonitor_66_or186;
  assign TLMonitor_66_or45 = TLMonitor_66_or91 | TLMonitor_66_or92;
  assign TLMonitor_66_or188 = stopEn83 | stopEn84;
  assign TLMonitor_66_or93 = stopEn82 | TLMonitor_66_or188;
  assign TLMonitor_66_or190 = stopEn86 | stopEn87;
  assign TLMonitor_66_or94 = stopEn85 | TLMonitor_66_or190;
  assign TLMonitor_66_or46 = TLMonitor_66_or93 | TLMonitor_66_or94;
  assign TLMonitor_66_or22 = TLMonitor_66_or45 | TLMonitor_66_or46;
  assign TLMonitor_66_or10 = TLMonitor_66_or21 | TLMonitor_66_or22;
  assign TLMonitor_66_or4 = TLMonitor_66_or9 | TLMonitor_66_or10;
  assign TLMonitor_66_or1 = TLMonitor_66_or3 | TLMonitor_66_or4;
  assign TLMonitor_66_or95 = stopEn88 | stopEn89;
  assign TLMonitor_66_or194 = stopEn91 | stopEn92;
  assign TLMonitor_66_or96 = stopEn90 | TLMonitor_66_or194;
  assign TLMonitor_66_or47 = TLMonitor_66_or95 | TLMonitor_66_or96;
  assign TLMonitor_66_or196 = stopEn94 | stopEn95;
  assign TLMonitor_66_or97 = stopEn93 | TLMonitor_66_or196;
  assign TLMonitor_66_or198 = stopEn97 | stopEn98;
  assign TLMonitor_66_or98 = stopEn96 | TLMonitor_66_or198;
  assign TLMonitor_66_or48 = TLMonitor_66_or97 | TLMonitor_66_or98;
  assign TLMonitor_66_or23 = TLMonitor_66_or47 | TLMonitor_66_or48;
  assign TLMonitor_66_or99 = stopEn99 | stopEn100;
  assign TLMonitor_66_or202 = stopEn102 | stopEn103;
  assign TLMonitor_66_or100 = stopEn101 | TLMonitor_66_or202;
  assign TLMonitor_66_or49 = TLMonitor_66_or99 | TLMonitor_66_or100;
  assign TLMonitor_66_or204 = stopEn105 | stopEn106;
  assign TLMonitor_66_or101 = stopEn104 | TLMonitor_66_or204;
  assign TLMonitor_66_or206 = stopEn108 | stopEn109;
  assign TLMonitor_66_or102 = stopEn107 | TLMonitor_66_or206;
  assign TLMonitor_66_or50 = TLMonitor_66_or101 | TLMonitor_66_or102;
  assign TLMonitor_66_or24 = TLMonitor_66_or49 | TLMonitor_66_or50;
  assign TLMonitor_66_or11 = TLMonitor_66_or23 | TLMonitor_66_or24;
  assign TLMonitor_66_or103 = stopEn110 | stopEn111;
  assign TLMonitor_66_or210 = stopEn113 | stopEn114;
  assign TLMonitor_66_or104 = stopEn112 | TLMonitor_66_or210;
  assign TLMonitor_66_or51 = TLMonitor_66_or103 | TLMonitor_66_or104;
  assign TLMonitor_66_or212 = stopEn116 | stopEn117;
  assign TLMonitor_66_or105 = stopEn115 | TLMonitor_66_or212;
  assign TLMonitor_66_or214 = stopEn119 | stopEn120;
  assign TLMonitor_66_or106 = stopEn118 | TLMonitor_66_or214;
  assign TLMonitor_66_or52 = TLMonitor_66_or105 | TLMonitor_66_or106;
  assign TLMonitor_66_or25 = TLMonitor_66_or51 | TLMonitor_66_or52;
  assign TLMonitor_66_or107 = stopEn121 | stopEn122;
  assign TLMonitor_66_or218 = stopEn124 | stopEn125;
  assign TLMonitor_66_or108 = stopEn123 | TLMonitor_66_or218;
  assign TLMonitor_66_or53 = TLMonitor_66_or107 | TLMonitor_66_or108;
  assign TLMonitor_66_or220 = stopEn127 | stopEn128;
  assign TLMonitor_66_or109 = stopEn126 | TLMonitor_66_or220;
  assign TLMonitor_66_or222 = stopEn130 | stopEn131;
  assign TLMonitor_66_or110 = stopEn129 | TLMonitor_66_or222;
  assign TLMonitor_66_or54 = TLMonitor_66_or109 | TLMonitor_66_or110;
  assign TLMonitor_66_or26 = TLMonitor_66_or53 | TLMonitor_66_or54;
  assign TLMonitor_66_or12 = TLMonitor_66_or25 | TLMonitor_66_or26;
  assign TLMonitor_66_or5 = TLMonitor_66_or11 | TLMonitor_66_or12;
  assign TLMonitor_66_or111 = stopEn132 | stopEn133;
  assign TLMonitor_66_or226 = stopEn135 | stopEn136;
  assign TLMonitor_66_or112 = stopEn134 | TLMonitor_66_or226;
  assign TLMonitor_66_or55 = TLMonitor_66_or111 | TLMonitor_66_or112;
  assign TLMonitor_66_or228 = stopEn138 | stopEn139;
  assign TLMonitor_66_or113 = stopEn137 | TLMonitor_66_or228;
  assign TLMonitor_66_or230 = stopEn141 | stopEn142;
  assign TLMonitor_66_or114 = stopEn140 | TLMonitor_66_or230;
  assign TLMonitor_66_or56 = TLMonitor_66_or113 | TLMonitor_66_or114;
  assign TLMonitor_66_or27 = TLMonitor_66_or55 | TLMonitor_66_or56;
  assign TLMonitor_66_or115 = stopEn143 | stopEn144;
  assign TLMonitor_66_or234 = stopEn146 | stopEn147;
  assign TLMonitor_66_or116 = stopEn145 | TLMonitor_66_or234;
  assign TLMonitor_66_or57 = TLMonitor_66_or115 | TLMonitor_66_or116;
  assign TLMonitor_66_or236 = stopEn149 | stopEn150;
  assign TLMonitor_66_or117 = stopEn148 | TLMonitor_66_or236;
  assign TLMonitor_66_or238 = stopEn152 | stopEn153;
  assign TLMonitor_66_or118 = stopEn151 | TLMonitor_66_or238;
  assign TLMonitor_66_or58 = TLMonitor_66_or117 | TLMonitor_66_or118;
  assign TLMonitor_66_or28 = TLMonitor_66_or57 | TLMonitor_66_or58;
  assign TLMonitor_66_or13 = TLMonitor_66_or27 | TLMonitor_66_or28;
  assign TLMonitor_66_or119 = stopEn154 | stopEn155;
  assign TLMonitor_66_or242 = stopEn157 | stopEn158;
  assign TLMonitor_66_or120 = stopEn156 | TLMonitor_66_or242;
  assign TLMonitor_66_or59 = TLMonitor_66_or119 | TLMonitor_66_or120;
  assign TLMonitor_66_or244 = stopEn160 | stopEn161;
  assign TLMonitor_66_or121 = stopEn159 | TLMonitor_66_or244;
  assign TLMonitor_66_or246 = stopEn163 | stopEn164;
  assign TLMonitor_66_or122 = stopEn162 | TLMonitor_66_or246;
  assign TLMonitor_66_or60 = TLMonitor_66_or121 | TLMonitor_66_or122;
  assign TLMonitor_66_or29 = TLMonitor_66_or59 | TLMonitor_66_or60;
  assign TLMonitor_66_or123 = stopEn165 | stopEn166;
  assign TLMonitor_66_or250 = stopEn168 | stopEn169;
  assign TLMonitor_66_or124 = stopEn167 | TLMonitor_66_or250;
  assign TLMonitor_66_or61 = TLMonitor_66_or123 | TLMonitor_66_or124;
  assign TLMonitor_66_or252 = stopEn171 | stopEn172;
  assign TLMonitor_66_or125 = stopEn170 | TLMonitor_66_or252;
  assign TLMonitor_66_or254 = stopEn174 | stopEn175;
  assign TLMonitor_66_or126 = stopEn173 | TLMonitor_66_or254;
  assign TLMonitor_66_or62 = TLMonitor_66_or125 | TLMonitor_66_or126;
  assign TLMonitor_66_or30 = TLMonitor_66_or61 | TLMonitor_66_or62;
  assign TLMonitor_66_or14 = TLMonitor_66_or29 | TLMonitor_66_or30;
  assign TLMonitor_66_or6 = TLMonitor_66_or13 | TLMonitor_66_or14;
  assign TLMonitor_66_or2 = TLMonitor_66_or5 | TLMonitor_66_or6;
  assign TLMonitor_66_or0 = TLMonitor_66_or1 | TLMonitor_66_or2;
  assign metaAssert = TLMonitor_66_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1669 = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1682 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1684 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1686 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1688 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1690 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_1724 = _RAND_6[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_1737 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_1739 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_1741 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_1743 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_1745 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_1747 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_1786 = _RAND_13[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_1799 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_1801 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_1803 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_1805 = _RAND_17[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_1807 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_1841 = _RAND_19[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_1854 = _RAND_20[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_1856 = _RAND_21[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_1858 = _RAND_22[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_1860 = _RAND_23[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_1862 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_1888 = _RAND_25[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_1899 = _RAND_26[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_1920 = _RAND_27[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_1986 = _RAND_28[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_1996 = _RAND_29[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  TLMonitor_66_metaAssert = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      _T_1669 <= 9'h0;
    end else if (reset) begin
      _T_1669 <= 9'h0;
    end else if (_T_1659) begin
      if (_T_1673) begin
        if (~io_in_a_bits_opcode[2]) begin
          _T_1669 <= _T_1664;
        end else begin
          _T_1669 <= 9'h0;
        end
      end else begin
        _T_1669 <= _T_1672;
      end
    end
    if (metaReset) begin
      _T_1682 <= 3'h0;
    end else if (_T_1714) begin
      _T_1682 <= io_in_a_bits_opcode;
    end
    if (metaReset) begin
      _T_1684 <= 3'h0;
    end else if (_T_1714) begin
      _T_1684 <= io_in_a_bits_param;
    end
    if (metaReset) begin
      _T_1686 <= 4'h0;
    end else if (_T_1714) begin
      _T_1686 <= io_in_a_bits_size;
    end
    if (metaReset) begin
      _T_1688 <= 2'h0;
    end else if (_T_1714) begin
      _T_1688 <= io_in_a_bits_source;
    end
    if (metaReset) begin
      _T_1690 <= 32'h0;
    end else if (_T_1714) begin
      _T_1690 <= io_in_a_bits_address;
    end
    if (metaReset) begin
      _T_1724 <= 9'h0;
    end else if (reset) begin
      _T_1724 <= 9'h0;
    end else if (_T_1715) begin
      if (_T_1728) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1724 <= _T_1720;
        end else begin
          _T_1724 <= 9'h0;
        end
      end else begin
        _T_1724 <= _T_1727;
      end
    end
    if (metaReset) begin
      _T_1737 <= 3'h0;
    end else if (_T_1775) begin
      _T_1737 <= io_in_d_bits_opcode;
    end
    if (metaReset) begin
      _T_1739 <= 2'h0;
    end else if (_T_1775) begin
      _T_1739 <= io_in_d_bits_param;
    end
    if (metaReset) begin
      _T_1741 <= 4'h0;
    end else if (_T_1775) begin
      _T_1741 <= io_in_d_bits_size;
    end
    if (metaReset) begin
      _T_1743 <= 2'h0;
    end else if (_T_1775) begin
      _T_1743 <= io_in_d_bits_source;
    end
    if (metaReset) begin
      _T_1745 <= 2'h0;
    end else if (_T_1775) begin
      _T_1745 <= io_in_d_bits_sink;
    end
    if (metaReset) begin
      _T_1747 <= 1'h0;
    end else if (_T_1775) begin
      _T_1747 <= io_in_d_bits_denied;
    end
    if (metaReset) begin
      _T_1786 <= 9'h0;
    end else if (reset) begin
      _T_1786 <= 9'h0;
    end else if (_T_1776) begin
      if (_T_1790) begin
        _T_1786 <= 9'h0;
      end else begin
        _T_1786 <= _T_1789;
      end
    end
    if (metaReset) begin
      _T_1799 <= 3'h0;
    end else if (_T_1831) begin
      _T_1799 <= io_in_b_bits_opcode;
    end
    if (metaReset) begin
      _T_1801 <= 2'h0;
    end else if (_T_1831) begin
      _T_1801 <= io_in_b_bits_param;
    end
    if (metaReset) begin
      _T_1803 <= 4'h0;
    end else if (_T_1831) begin
      _T_1803 <= io_in_b_bits_size;
    end
    if (metaReset) begin
      _T_1805 <= 2'h0;
    end else if (_T_1831) begin
      _T_1805 <= io_in_b_bits_source;
    end
    if (metaReset) begin
      _T_1807 <= 32'h0;
    end else if (_T_1831) begin
      _T_1807 <= io_in_b_bits_address;
    end
    if (metaReset) begin
      _T_1841 <= 9'h0;
    end else if (reset) begin
      _T_1841 <= 9'h0;
    end else if (_T_1832) begin
      if (_T_1845) begin
        if (io_in_c_bits_opcode[0]) begin
          _T_1841 <= _T_1837;
        end else begin
          _T_1841 <= 9'h0;
        end
      end else begin
        _T_1841 <= _T_1844;
      end
    end
    if (metaReset) begin
      _T_1854 <= 3'h0;
    end else if (_T_1886) begin
      _T_1854 <= io_in_c_bits_opcode;
    end
    if (metaReset) begin
      _T_1856 <= 3'h0;
    end else if (_T_1886) begin
      _T_1856 <= io_in_c_bits_param;
    end
    if (metaReset) begin
      _T_1858 <= 4'h0;
    end else if (_T_1886) begin
      _T_1858 <= io_in_c_bits_size;
    end
    if (metaReset) begin
      _T_1860 <= 2'h0;
    end else if (_T_1886) begin
      _T_1860 <= io_in_c_bits_source;
    end
    if (metaReset) begin
      _T_1862 <= 32'h0;
    end else if (_T_1886) begin
      _T_1862 <= io_in_c_bits_address;
    end
    if (metaReset) begin
      _T_1888 <= 3'h0;
    end else if (reset) begin
      _T_1888 <= 3'h0;
    end else begin
      _T_1888 <= _T_1968;
    end
    if (metaReset) begin
      _T_1899 <= 9'h0;
    end else if (reset) begin
      _T_1899 <= 9'h0;
    end else if (_T_1659) begin
      if (_T_1903) begin
        if (~io_in_a_bits_opcode[2]) begin
          _T_1899 <= _T_1664;
        end else begin
          _T_1899 <= 9'h0;
        end
      end else begin
        _T_1899 <= _T_1902;
      end
    end
    if (metaReset) begin
      _T_1920 <= 9'h0;
    end else if (reset) begin
      _T_1920 <= 9'h0;
    end else if (_T_1715) begin
      if (_T_1924) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1920 <= _T_1720;
        end else begin
          _T_1920 <= 9'h0;
        end
      end else begin
        _T_1920 <= _T_1923;
      end
    end
    if (metaReset) begin
      _T_1986 <= 4'h0;
    end else if (reset) begin
      _T_1986 <= 4'h0;
    end else begin
      _T_1986 <= _T_2038;
    end
    if (metaReset) begin
      _T_1996 <= 9'h0;
    end else if (reset) begin
      _T_1996 <= 9'h0;
    end else if (_T_1715) begin
      if (_T_2000) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1996 <= _T_1720;
        end else begin
          _T_1996 <= 9'h0;
        end
      end else begin
        _T_1996 <= _T_1999;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_37 & ~_T_184) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:49 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquireBlock type unsupported by manager\" + extra)\n"); // @[Monitor.scala 49:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_37 & ~_T_184) begin
          $fatal; // @[Monitor.scala 49:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_37 & ~_T_208) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:50 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquireBlock from a client which does not support Probe\" + extra)\n"); // @[Monitor.scala 50:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_37 & ~_T_208) begin
          $fatal; // @[Monitor.scala 50:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_37 & ~_T_211) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert (source_ok, \"'A' channel AcquireBlock carries invalid source ID\" + extra)\n"); // @[Monitor.scala 51:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_37 & ~_T_211) begin
          $fatal; // @[Monitor.scala 51:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_37 & ~_T_215) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:52 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquireBlock smaller than a beat\" + extra)\n"); // @[Monitor.scala 52:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_37 & ~_T_215) begin
          $fatal; // @[Monitor.scala 52:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_37 & ~_T_218) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:53 assert (is_aligned, \"'A' channel AcquireBlock address not aligned to size\" + extra)\n"); // @[Monitor.scala 53:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_37 & ~_T_218) begin
          $fatal; // @[Monitor.scala 53:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_37 & ~_T_222) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:54 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquireBlock carries invalid grow param\" + extra)\n"); // @[Monitor.scala 54:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_37 & ~_T_222) begin
          $fatal; // @[Monitor.scala 54:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_37 & ~_T_227) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:55 assert (~bundle.mask === UInt(0), \"'A' channel AcquireBlock contains invalid mask\" + extra)\n"); // @[Monitor.scala 55:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_37 & ~_T_227) begin
          $fatal; // @[Monitor.scala 55:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_37 & ~_T_231) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:56 assert (!bundle.corrupt, \"'A' channel AcquireBlock is corrupt\" + extra)\n"); // @[Monitor.scala 56:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_37 & ~_T_231) begin
          $fatal; // @[Monitor.scala 56:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & ~_T_184) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:60 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquirePerm type unsupported by manager\" + extra)\n"); // @[Monitor.scala 60:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & ~_T_184) begin
          $fatal; // @[Monitor.scala 60:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & ~_T_208) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:61 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquirePerm from a client which does not support Probe\" + extra)\n"); // @[Monitor.scala 61:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & ~_T_208) begin
          $fatal; // @[Monitor.scala 61:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & ~_T_211) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:62 assert (source_ok, \"'A' channel AcquirePerm carries invalid source ID\" + extra)\n"); // @[Monitor.scala 62:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & ~_T_211) begin
          $fatal; // @[Monitor.scala 62:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & ~_T_215) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:63 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquirePerm smaller than a beat\" + extra)\n"); // @[Monitor.scala 63:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & ~_T_215) begin
          $fatal; // @[Monitor.scala 63:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & ~_T_218) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:64 assert (is_aligned, \"'A' channel AcquirePerm address not aligned to size\" + extra)\n"); // @[Monitor.scala 64:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & ~_T_218) begin
          $fatal; // @[Monitor.scala 64:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & ~_T_222) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:65 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquirePerm carries invalid grow param\" + extra)\n"); // @[Monitor.scala 65:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & ~_T_222) begin
          $fatal; // @[Monitor.scala 65:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & ~_T_326) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:66 assert (bundle.param =/= TLPermissions.NtoB, \"'A' channel AcquirePerm requests NtoB\" + extra)\n"); // @[Monitor.scala 66:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & ~_T_326) begin
          $fatal; // @[Monitor.scala 66:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & ~_T_227) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:67 assert (~bundle.mask === UInt(0), \"'A' channel AcquirePerm contains invalid mask\" + extra)\n"); // @[Monitor.scala 67:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & ~_T_227) begin
          $fatal; // @[Monitor.scala 67:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & ~_T_231) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:68 assert (!bundle.corrupt, \"'A' channel AcquirePerm is corrupt\" + extra)\n"); // @[Monitor.scala 68:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & ~_T_231) begin
          $fatal; // @[Monitor.scala 68:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_71 & ~_T_391) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:72 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); // @[Monitor.scala 72:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_71 & ~_T_391) begin
          $fatal; // @[Monitor.scala 72:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_71 & ~_T_211) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:73 assert (source_ok, \"'A' channel Get carries invalid source ID\" + extra)\n"); // @[Monitor.scala 73:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_71 & ~_T_211) begin
          $fatal; // @[Monitor.scala 73:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_71 & ~_T_218) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:74 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); // @[Monitor.scala 74:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_71 & ~_T_218) begin
          $fatal; // @[Monitor.scala 74:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_71 & ~_T_401) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:75 assert (bundle.param === UInt(0), \"'A' channel Get carries invalid param\" + extra)\n"); // @[Monitor.scala 75:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_71 & ~_T_401) begin
          $fatal; // @[Monitor.scala 75:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_71 & ~_T_405) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:76 assert (bundle.mask === mask, \"'A' channel Get contains invalid mask\" + extra)\n"); // @[Monitor.scala 76:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_71 & ~_T_405) begin
          $fatal; // @[Monitor.scala 76:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_71 & ~_T_231) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:77 assert (!bundle.corrupt, \"'A' channel Get is corrupt\" + extra)\n"); // @[Monitor.scala 77:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_71 & ~_T_231) begin
          $fatal; // @[Monitor.scala 77:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_83 & ~_T_472) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:81 assert (edge.manager.supportsPutFullSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutFull type unsupported by manager\" + extra)\n"); // @[Monitor.scala 81:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_83 & ~_T_472) begin
          $fatal; // @[Monitor.scala 81:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_83 & ~_T_211) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:82 assert (source_ok, \"'A' channel PutFull carries invalid source ID\" + extra)\n"); // @[Monitor.scala 82:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_83 & ~_T_211) begin
          $fatal; // @[Monitor.scala 82:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_83 & ~_T_218) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:83 assert (is_aligned, \"'A' channel PutFull address not aligned to size\" + extra)\n"); // @[Monitor.scala 83:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_83 & ~_T_218) begin
          $fatal; // @[Monitor.scala 83:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_83 & ~_T_401) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:84 assert (bundle.param === UInt(0), \"'A' channel PutFull carries invalid param\" + extra)\n"); // @[Monitor.scala 84:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_83 & ~_T_401) begin
          $fatal; // @[Monitor.scala 84:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_83 & ~_T_405) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:85 assert (bundle.mask === mask, \"'A' channel PutFull contains invalid mask\" + extra)\n"); // @[Monitor.scala 85:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_83 & ~_T_405) begin
          $fatal; // @[Monitor.scala 85:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & ~_T_472) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:89 assert (edge.manager.supportsPutPartialSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutPartial type unsupported by manager\" + extra)\n"); // @[Monitor.scala 89:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & ~_T_472) begin
          $fatal; // @[Monitor.scala 89:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & ~_T_211) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:90 assert (source_ok, \"'A' channel PutPartial carries invalid source ID\" + extra)\n"); // @[Monitor.scala 90:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & ~_T_211) begin
          $fatal; // @[Monitor.scala 90:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & ~_T_218) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:91 assert (is_aligned, \"'A' channel PutPartial address not aligned to size\" + extra)\n"); // @[Monitor.scala 91:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & ~_T_218) begin
          $fatal; // @[Monitor.scala 91:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & ~_T_401) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:92 assert (bundle.param === UInt(0), \"'A' channel PutPartial carries invalid param\" + extra)\n"); // @[Monitor.scala 92:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & ~_T_401) begin
          $fatal; // @[Monitor.scala 92:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & ~_T_565) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:93 assert ((bundle.mask & ~mask) === UInt(0), \"'A' channel PutPartial contains invalid mask\" + extra)\n"); // @[Monitor.scala 93:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & ~_T_565) begin
          $fatal; // @[Monitor.scala 93:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & ~_T_618) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:97 assert (edge.manager.supportsArithmeticSafe(edge.address(bundle), bundle.size), \"'A' channel carries Arithmetic type unsupported by manager\" + extra)\n"); // @[Monitor.scala 97:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & ~_T_618) begin
          $fatal; // @[Monitor.scala 97:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & ~_T_211) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:98 assert (source_ok, \"'A' channel Arithmetic carries invalid source ID\" + extra)\n"); // @[Monitor.scala 98:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & ~_T_211) begin
          $fatal; // @[Monitor.scala 98:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & ~_T_218) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:99 assert (is_aligned, \"'A' channel Arithmetic address not aligned to size\" + extra)\n"); // @[Monitor.scala 99:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & ~_T_218) begin
          $fatal; // @[Monitor.scala 99:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & ~_T_628) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:100 assert (TLAtomics.isArithmetic(bundle.param), \"'A' channel Arithmetic carries invalid opcode param\" + extra)\n"); // @[Monitor.scala 100:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & ~_T_628) begin
          $fatal; // @[Monitor.scala 100:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & ~_T_405) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:101 assert (bundle.mask === mask, \"'A' channel Arithmetic contains invalid mask\" + extra)\n"); // @[Monitor.scala 101:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & ~_T_405) begin
          $fatal; // @[Monitor.scala 101:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_113 & ~_T_618) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:105 assert (edge.manager.supportsLogicalSafe(edge.address(bundle), bundle.size), \"'A' channel carries Logical type unsupported by manager\" + extra)\n"); // @[Monitor.scala 105:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_113 & ~_T_618) begin
          $fatal; // @[Monitor.scala 105:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_113 & ~_T_211) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:106 assert (source_ok, \"'A' channel Logical carries invalid source ID\" + extra)\n"); // @[Monitor.scala 106:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_113 & ~_T_211) begin
          $fatal; // @[Monitor.scala 106:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_113 & ~_T_218) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:107 assert (is_aligned, \"'A' channel Logical address not aligned to size\" + extra)\n"); // @[Monitor.scala 107:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_113 & ~_T_218) begin
          $fatal; // @[Monitor.scala 107:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_113 & ~_T_695) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:108 assert (TLAtomics.isLogical(bundle.param), \"'A' channel Logical carries invalid opcode param\" + extra)\n"); // @[Monitor.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_113 & ~_T_695) begin
          $fatal; // @[Monitor.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_113 & ~_T_405) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:109 assert (bundle.mask === mask, \"'A' channel Logical contains invalid mask\" + extra)\n"); // @[Monitor.scala 109:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_113 & ~_T_405) begin
          $fatal; // @[Monitor.scala 109:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & ~_T_752) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:113 assert (edge.manager.supportsHintSafe(edge.address(bundle), bundle.size), \"'A' channel carries Hint type unsupported by manager\" + extra)\n"); // @[Monitor.scala 113:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & ~_T_752) begin
          $fatal; // @[Monitor.scala 113:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & ~_T_211) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:114 assert (source_ok, \"'A' channel Hint carries invalid source ID\" + extra)\n"); // @[Monitor.scala 114:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & ~_T_211) begin
          $fatal; // @[Monitor.scala 114:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & ~_T_218) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:115 assert (is_aligned, \"'A' channel Hint address not aligned to size\" + extra)\n"); // @[Monitor.scala 115:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & ~_T_218) begin
          $fatal; // @[Monitor.scala 115:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & ~_T_405) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:116 assert (bundle.mask === mask, \"'A' channel Hint contains invalid mask\" + extra)\n"); // @[Monitor.scala 116:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & ~_T_405) begin
          $fatal; // @[Monitor.scala 116:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & ~_T_231) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:117 assert (!bundle.corrupt, \"'A' channel Hint is corrupt\" + extra)\n"); // @[Monitor.scala 117:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & ~_T_231) begin
          $fatal; // @[Monitor.scala 117:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~_T_770) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:268 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); // @[Monitor.scala 268:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~_T_770) begin
          $fatal; // @[Monitor.scala 268:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & ~_T_789) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:276 assert (source_ok, \"'D' channel ReleaseAck carries invalid source ID\" + extra)\n"); // @[Monitor.scala 276:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & ~_T_789) begin
          $fatal; // @[Monitor.scala 276:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & ~_T_793) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:277 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); // @[Monitor.scala 277:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & ~_T_793) begin
          $fatal; // @[Monitor.scala 277:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & ~_T_797) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:278 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); // @[Monitor.scala 278:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & ~_T_797) begin
          $fatal; // @[Monitor.scala 278:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & ~_T_801) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:279 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); // @[Monitor.scala 279:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & ~_T_801) begin
          $fatal; // @[Monitor.scala 279:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & ~_T_805) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:280 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); // @[Monitor.scala 280:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & ~_T_805) begin
          $fatal; // @[Monitor.scala 280:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & ~_T_789) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:284 assert (source_ok, \"'D' channel Grant carries invalid source ID\" + extra)\n"); // @[Monitor.scala 284:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & ~_T_789) begin
          $fatal; // @[Monitor.scala 284:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & ~_T_793) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:286 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); // @[Monitor.scala 286:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & ~_T_793) begin
          $fatal; // @[Monitor.scala 286:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & ~_T_820) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:287 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); // @[Monitor.scala 287:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & ~_T_820) begin
          $fatal; // @[Monitor.scala 287:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & ~_T_824) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:288 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); // @[Monitor.scala 288:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & ~_T_824) begin
          $fatal; // @[Monitor.scala 288:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & ~_T_801) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:289 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); // @[Monitor.scala 289:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & ~_T_801) begin
          $fatal; // @[Monitor.scala 289:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & ~_T_789) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:294 assert (source_ok, \"'D' channel GrantData carries invalid source ID\" + extra)\n"); // @[Monitor.scala 294:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & ~_T_789) begin
          $fatal; // @[Monitor.scala 294:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & ~_T_793) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:296 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); // @[Monitor.scala 296:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & ~_T_793) begin
          $fatal; // @[Monitor.scala 296:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & ~_T_820) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:297 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); // @[Monitor.scala 297:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & ~_T_820) begin
          $fatal; // @[Monitor.scala 297:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & ~_T_824) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:298 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); // @[Monitor.scala 298:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & ~_T_824) begin
          $fatal; // @[Monitor.scala 298:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & ~_T_857) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:299 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); // @[Monitor.scala 299:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & ~_T_857) begin
          $fatal; // @[Monitor.scala 299:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & ~_T_789) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:304 assert (source_ok, \"'D' channel AccessAck carries invalid source ID\" + extra)\n"); // @[Monitor.scala 304:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & ~_T_789) begin
          $fatal; // @[Monitor.scala 304:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & ~_T_797) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:306 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); // @[Monitor.scala 306:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & ~_T_797) begin
          $fatal; // @[Monitor.scala 306:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & ~_T_801) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:307 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); // @[Monitor.scala 307:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & ~_T_801) begin
          $fatal; // @[Monitor.scala 307:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_169 & ~_T_789) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:312 assert (source_ok, \"'D' channel AccessAckData carries invalid source ID\" + extra)\n"); // @[Monitor.scala 312:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_169 & ~_T_789) begin
          $fatal; // @[Monitor.scala 312:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_169 & ~_T_797) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:314 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); // @[Monitor.scala 314:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_169 & ~_T_797) begin
          $fatal; // @[Monitor.scala 314:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_169 & ~_T_857) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:315 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); // @[Monitor.scala 315:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_169 & ~_T_857) begin
          $fatal; // @[Monitor.scala 315:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & ~_T_789) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:320 assert (source_ok, \"'D' channel HintAck carries invalid source ID\" + extra)\n"); // @[Monitor.scala 320:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & ~_T_789) begin
          $fatal; // @[Monitor.scala 320:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & ~_T_797) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:322 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); // @[Monitor.scala 322:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & ~_T_797) begin
          $fatal; // @[Monitor.scala 322:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & ~_T_801) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:323 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); // @[Monitor.scala 323:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & ~_T_801) begin
          $fatal; // @[Monitor.scala 323:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_b_valid & ~_T_918) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel has invalid opcode (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:122 assert (TLMessages.isB(bundle.opcode), \"'B' channel has invalid opcode\" + extra)\n"); // @[Monitor.scala 122:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_b_valid & ~_T_918) begin
          $fatal; // @[Monitor.scala 122:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & ~_T_1117) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Probe type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:133 assert (edge.client.supportsProbe(bundle.source, bundle.size), \"'B' channel carries Probe type unsupported by client\" + extra)\n"); // @[Monitor.scala 133:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & ~_T_1117) begin
          $fatal; // @[Monitor.scala 133:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & ~_T_1120) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:134 assert (address_ok, \"'B' channel Probe carries unmanaged address\" + extra)\n"); // @[Monitor.scala 134:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & ~_T_1120) begin
          $fatal; // @[Monitor.scala 134:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & ~_T_1123) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:135 assert (legal_source, \"'B' channel Probe carries source that is not first source\" + extra)\n"); // @[Monitor.scala 135:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & ~_T_1123) begin
          $fatal; // @[Monitor.scala 135:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & ~_T_1126) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:136 assert (is_aligned, \"'B' channel Probe address not aligned to size\" + extra)\n"); // @[Monitor.scala 136:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & ~_T_1126) begin
          $fatal; // @[Monitor.scala 136:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & ~_T_1130) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries invalid cap param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:137 assert (TLPermissions.isCap(bundle.param), \"'B' channel Probe carries invalid cap param\" + extra)\n"); // @[Monitor.scala 137:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & ~_T_1130) begin
          $fatal; // @[Monitor.scala 137:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & ~_T_1134) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:138 assert (bundle.mask === mask, \"'B' channel Probe contains invalid mask\" + extra)\n"); // @[Monitor.scala 138:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & ~_T_1134) begin
          $fatal; // @[Monitor.scala 138:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & ~_T_1138) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:139 assert (!bundle.corrupt, \"'B' channel Probe is corrupt\" + extra)\n"); // @[Monitor.scala 139:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & ~_T_1138) begin
          $fatal; // @[Monitor.scala 139:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Get type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:143 assert (edge.client.supportsGet(bundle.source, bundle.size), \"'B' channel carries Get type unsupported by client\" + extra)\n"); // @[Monitor.scala 143:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & ~reset) begin
          $fatal; // @[Monitor.scala 143:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & ~_T_1120) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:144 assert (address_ok, \"'B' channel Get carries unmanaged address\" + extra)\n"); // @[Monitor.scala 144:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & ~_T_1120) begin
          $fatal; // @[Monitor.scala 144:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & ~_T_1123) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:145 assert (legal_source, \"'B' channel Get carries source that is not first source\" + extra)\n"); // @[Monitor.scala 145:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & ~_T_1123) begin
          $fatal; // @[Monitor.scala 145:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & ~_T_1126) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:146 assert (is_aligned, \"'B' channel Get address not aligned to size\" + extra)\n"); // @[Monitor.scala 146:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & ~_T_1126) begin
          $fatal; // @[Monitor.scala 146:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & ~_T_1155) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:147 assert (bundle.param === UInt(0), \"'B' channel Get carries invalid param\" + extra)\n"); // @[Monitor.scala 147:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & ~_T_1155) begin
          $fatal; // @[Monitor.scala 147:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & ~_T_1134) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:148 assert (bundle.mask === mask, \"'B' channel Get contains invalid mask\" + extra)\n"); // @[Monitor.scala 148:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & ~_T_1134) begin
          $fatal; // @[Monitor.scala 148:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & ~_T_1138) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:149 assert (!bundle.corrupt, \"'B' channel Get is corrupt\" + extra)\n"); // @[Monitor.scala 149:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & ~_T_1138) begin
          $fatal; // @[Monitor.scala 149:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_209 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutFull type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:153 assert (edge.client.supportsPutFull(bundle.source, bundle.size), \"'B' channel carries PutFull type unsupported by client\" + extra)\n"); // @[Monitor.scala 153:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_209 & ~reset) begin
          $fatal; // @[Monitor.scala 153:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_209 & ~_T_1120) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:154 assert (address_ok, \"'B' channel PutFull carries unmanaged address\" + extra)\n"); // @[Monitor.scala 154:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_209 & ~_T_1120) begin
          $fatal; // @[Monitor.scala 154:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_209 & ~_T_1123) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:155 assert (legal_source, \"'B' channel PutFull carries source that is not first source\" + extra)\n"); // @[Monitor.scala 155:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_209 & ~_T_1123) begin
          $fatal; // @[Monitor.scala 155:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_209 & ~_T_1126) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:156 assert (is_aligned, \"'B' channel PutFull address not aligned to size\" + extra)\n"); // @[Monitor.scala 156:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_209 & ~_T_1126) begin
          $fatal; // @[Monitor.scala 156:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_209 & ~_T_1155) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:157 assert (bundle.param === UInt(0), \"'B' channel PutFull carries invalid param\" + extra)\n"); // @[Monitor.scala 157:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_209 & ~_T_1155) begin
          $fatal; // @[Monitor.scala 157:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_209 & ~_T_1134) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:158 assert (bundle.mask === mask, \"'B' channel PutFull contains invalid mask\" + extra)\n"); // @[Monitor.scala 158:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_209 & ~_T_1134) begin
          $fatal; // @[Monitor.scala 158:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_221 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutPartial type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:162 assert (edge.client.supportsPutPartial(bundle.source, bundle.size), \"'B' channel carries PutPartial type unsupported by client\" + extra)\n"); // @[Monitor.scala 162:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_221 & ~reset) begin
          $fatal; // @[Monitor.scala 162:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_221 & ~_T_1120) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:163 assert (address_ok, \"'B' channel PutPartial carries unmanaged address\" + extra)\n"); // @[Monitor.scala 163:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_221 & ~_T_1120) begin
          $fatal; // @[Monitor.scala 163:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_221 & ~_T_1123) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:164 assert (legal_source, \"'B' channel PutPartial carries source that is not first source\" + extra)\n"); // @[Monitor.scala 164:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_221 & ~_T_1123) begin
          $fatal; // @[Monitor.scala 164:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_221 & ~_T_1126) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:165 assert (is_aligned, \"'B' channel PutPartial address not aligned to size\" + extra)\n"); // @[Monitor.scala 165:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_221 & ~_T_1126) begin
          $fatal; // @[Monitor.scala 165:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_221 & ~_T_1155) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:166 assert (bundle.param === UInt(0), \"'B' channel PutPartial carries invalid param\" + extra)\n"); // @[Monitor.scala 166:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_221 & ~_T_1155) begin
          $fatal; // @[Monitor.scala 166:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_221 & ~_T_1207) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:167 assert ((bundle.mask & ~mask) === UInt(0), \"'B' channel PutPartial contains invalid mask\" + extra)\n"); // @[Monitor.scala 167:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_221 & ~_T_1207) begin
          $fatal; // @[Monitor.scala 167:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Arithmetic type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:171 assert (edge.client.supportsArithmetic(bundle.source, bundle.size), \"'B' channel carries Arithmetic type unsupported by client\" + extra)\n"); // @[Monitor.scala 171:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & ~reset) begin
          $fatal; // @[Monitor.scala 171:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & ~_T_1120) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:172 assert (address_ok, \"'B' channel Arithmetic carries unmanaged address\" + extra)\n"); // @[Monitor.scala 172:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & ~_T_1120) begin
          $fatal; // @[Monitor.scala 172:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & ~_T_1123) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:173 assert (legal_source, \"'B' channel Arithmetic carries source that is not first source\" + extra)\n"); // @[Monitor.scala 173:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & ~_T_1123) begin
          $fatal; // @[Monitor.scala 173:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & ~_T_1126) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:174 assert (is_aligned, \"'B' channel Arithmetic address not aligned to size\" + extra)\n"); // @[Monitor.scala 174:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & ~_T_1126) begin
          $fatal; // @[Monitor.scala 174:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & ~_T_1134) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:176 assert (bundle.mask === mask, \"'B' channel Arithmetic contains invalid mask\" + extra)\n"); // @[Monitor.scala 176:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & ~_T_1134) begin
          $fatal; // @[Monitor.scala 176:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_243 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Logical type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:180 assert (edge.client.supportsLogical(bundle.source, bundle.size), \"'B' channel carries Logical type unsupported by client\" + extra)\n"); // @[Monitor.scala 180:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_243 & ~reset) begin
          $fatal; // @[Monitor.scala 180:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_243 & ~_T_1120) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:181 assert (address_ok, \"'B' channel Logical carries unmanaged address\" + extra)\n"); // @[Monitor.scala 181:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_243 & ~_T_1120) begin
          $fatal; // @[Monitor.scala 181:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_243 & ~_T_1123) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:182 assert (legal_source, \"'B' channel Logical carries source that is not first source\" + extra)\n"); // @[Monitor.scala 182:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_243 & ~_T_1123) begin
          $fatal; // @[Monitor.scala 182:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_243 & ~_T_1126) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:183 assert (is_aligned, \"'B' channel Logical address not aligned to size\" + extra)\n"); // @[Monitor.scala 183:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_243 & ~_T_1126) begin
          $fatal; // @[Monitor.scala 183:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_243 & ~_T_1134) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:185 assert (bundle.mask === mask, \"'B' channel Logical contains invalid mask\" + extra)\n"); // @[Monitor.scala 185:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_243 & ~_T_1134) begin
          $fatal; // @[Monitor.scala 185:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_253 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Hint type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:189 assert (edge.client.supportsHint(bundle.source, bundle.size), \"'B' channel carries Hint type unsupported by client\" + extra)\n"); // @[Monitor.scala 189:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_253 & ~reset) begin
          $fatal; // @[Monitor.scala 189:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_253 & ~_T_1120) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:190 assert (address_ok, \"'B' channel Hint carries unmanaged address\" + extra)\n"); // @[Monitor.scala 190:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_253 & ~_T_1120) begin
          $fatal; // @[Monitor.scala 190:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_253 & ~_T_1123) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:191 assert (legal_source, \"'B' channel Hint carries source that is not first source\" + extra)\n"); // @[Monitor.scala 191:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_253 & ~_T_1123) begin
          $fatal; // @[Monitor.scala 191:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_253 & ~_T_1126) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:192 assert (is_aligned, \"'B' channel Hint address not aligned to size\" + extra)\n"); // @[Monitor.scala 192:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_253 & ~_T_1126) begin
          $fatal; // @[Monitor.scala 192:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_253 & ~_T_1134) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:193 assert (bundle.mask === mask, \"'B' channel Hint contains invalid mask\" + extra)\n"); // @[Monitor.scala 193:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_253 & ~_T_1134) begin
          $fatal; // @[Monitor.scala 193:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_253 & ~_T_1138) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:194 assert (!bundle.corrupt, \"'B' channel Hint is corrupt\" + extra)\n"); // @[Monitor.scala 194:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_253 & ~_T_1138) begin
          $fatal; // @[Monitor.scala 194:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_265 & ~_T_1381) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:208 assert (address_ok, \"'C' channel ProbeAck carries unmanaged address\" + extra)\n"); // @[Monitor.scala 208:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & ~_T_1381) begin
          $fatal; // @[Monitor.scala 208:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_265 & ~_T_1384) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:209 assert (source_ok, \"'C' channel ProbeAck carries invalid source ID\" + extra)\n"); // @[Monitor.scala 209:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & ~_T_1384) begin
          $fatal; // @[Monitor.scala 209:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_265 & ~_T_1388) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:210 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAck smaller than a beat\" + extra)\n"); // @[Monitor.scala 210:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & ~_T_1388) begin
          $fatal; // @[Monitor.scala 210:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_265 & ~_T_1391) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:211 assert (is_aligned, \"'C' channel ProbeAck address not aligned to size\" + extra)\n"); // @[Monitor.scala 211:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & ~_T_1391) begin
          $fatal; // @[Monitor.scala 211:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_265 & ~_T_1395) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:212 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAck carries invalid report param\" + extra)\n"); // @[Monitor.scala 212:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & ~_T_1395) begin
          $fatal; // @[Monitor.scala 212:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_275 & ~_T_1381) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:217 assert (address_ok, \"'C' channel ProbeAckData carries unmanaged address\" + extra)\n"); // @[Monitor.scala 217:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_275 & ~_T_1381) begin
          $fatal; // @[Monitor.scala 217:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_275 & ~_T_1384) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:218 assert (source_ok, \"'C' channel ProbeAckData carries invalid source ID\" + extra)\n"); // @[Monitor.scala 218:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_275 & ~_T_1384) begin
          $fatal; // @[Monitor.scala 218:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_275 & ~_T_1388) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:219 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAckData smaller than a beat\" + extra)\n"); // @[Monitor.scala 219:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_275 & ~_T_1388) begin
          $fatal; // @[Monitor.scala 219:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_275 & ~_T_1391) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:220 assert (is_aligned, \"'C' channel ProbeAckData address not aligned to size\" + extra)\n"); // @[Monitor.scala 220:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_275 & ~_T_1391) begin
          $fatal; // @[Monitor.scala 220:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_275 & ~_T_1395) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:221 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAckData carries invalid report param\" + extra)\n"); // @[Monitor.scala 221:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_275 & ~_T_1395) begin
          $fatal; // @[Monitor.scala 221:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & ~_T_1470) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:225 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries Release type unsupported by manager\" + extra)\n"); // @[Monitor.scala 225:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & ~_T_1470) begin
          $fatal; // @[Monitor.scala 225:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & ~_T_1494) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:226 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); // @[Monitor.scala 226:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & ~_T_1494) begin
          $fatal; // @[Monitor.scala 226:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & ~_T_1384) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:227 assert (source_ok, \"'C' channel Release carries invalid source ID\" + extra)\n"); // @[Monitor.scala 227:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & ~_T_1384) begin
          $fatal; // @[Monitor.scala 227:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & ~_T_1388) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:228 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel Release smaller than a beat\" + extra)\n"); // @[Monitor.scala 228:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & ~_T_1388) begin
          $fatal; // @[Monitor.scala 228:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & ~_T_1391) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:229 assert (is_aligned, \"'C' channel Release address not aligned to size\" + extra)\n"); // @[Monitor.scala 229:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & ~_T_1391) begin
          $fatal; // @[Monitor.scala 229:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & ~_T_1508) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid shrink param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:230 assert (TLPermissions.isShrink(bundle.param), \"'C' channel Release carries invalid shrink param\" + extra)\n"); // @[Monitor.scala 230:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & ~_T_1508) begin
          $fatal; // @[Monitor.scala 230:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_297 & ~_T_1470) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:235 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries ReleaseData type unsupported by manager\" + extra)\n"); // @[Monitor.scala 235:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_297 & ~_T_1470) begin
          $fatal; // @[Monitor.scala 235:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_297 & ~_T_1494) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:236 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); // @[Monitor.scala 236:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_297 & ~_T_1494) begin
          $fatal; // @[Monitor.scala 236:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_297 & ~_T_1384) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:237 assert (source_ok, \"'C' channel ReleaseData carries invalid source ID\" + extra)\n"); // @[Monitor.scala 237:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_297 & ~_T_1384) begin
          $fatal; // @[Monitor.scala 237:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_297 & ~_T_1388) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:238 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ReleaseData smaller than a beat\" + extra)\n"); // @[Monitor.scala 238:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_297 & ~_T_1388) begin
          $fatal; // @[Monitor.scala 238:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_297 & ~_T_1391) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:239 assert (is_aligned, \"'C' channel ReleaseData address not aligned to size\" + extra)\n"); // @[Monitor.scala 239:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_297 & ~_T_1391) begin
          $fatal; // @[Monitor.scala 239:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_297 & ~_T_1508) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid shrink param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:240 assert (TLPermissions.isShrink(bundle.param), \"'C' channel ReleaseData carries invalid shrink param\" + extra)\n"); // @[Monitor.scala 240:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_297 & ~_T_1508) begin
          $fatal; // @[Monitor.scala 240:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_309 & ~_T_1381) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:244 assert (address_ok, \"'C' channel AccessAck carries unmanaged address\" + extra)\n"); // @[Monitor.scala 244:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_309 & ~_T_1381) begin
          $fatal; // @[Monitor.scala 244:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_309 & ~_T_1384) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:245 assert (source_ok, \"'C' channel AccessAck carries invalid source ID\" + extra)\n"); // @[Monitor.scala 245:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_309 & ~_T_1384) begin
          $fatal; // @[Monitor.scala 245:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_309 & ~_T_1391) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:246 assert (is_aligned, \"'C' channel AccessAck address not aligned to size\" + extra)\n"); // @[Monitor.scala 246:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_309 & ~_T_1391) begin
          $fatal; // @[Monitor.scala 246:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_309 & ~_T_1617) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:247 assert (bundle.param === UInt(0), \"'C' channel AccessAck carries invalid param\" + extra)\n"); // @[Monitor.scala 247:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_309 & ~_T_1617) begin
          $fatal; // @[Monitor.scala 247:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & ~_T_1381) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:252 assert (address_ok, \"'C' channel AccessAckData carries unmanaged address\" + extra)\n"); // @[Monitor.scala 252:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & ~_T_1381) begin
          $fatal; // @[Monitor.scala 252:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & ~_T_1384) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:253 assert (source_ok, \"'C' channel AccessAckData carries invalid source ID\" + extra)\n"); // @[Monitor.scala 253:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & ~_T_1384) begin
          $fatal; // @[Monitor.scala 253:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & ~_T_1391) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:254 assert (is_aligned, \"'C' channel AccessAckData address not aligned to size\" + extra)\n"); // @[Monitor.scala 254:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & ~_T_1391) begin
          $fatal; // @[Monitor.scala 254:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & ~_T_1617) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:255 assert (bundle.param === UInt(0), \"'C' channel AccessAckData carries invalid param\" + extra)\n"); // @[Monitor.scala 255:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & ~_T_1617) begin
          $fatal; // @[Monitor.scala 255:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_325 & ~_T_1381) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:259 assert (address_ok, \"'C' channel HintAck carries unmanaged address\" + extra)\n"); // @[Monitor.scala 259:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_325 & ~_T_1381) begin
          $fatal; // @[Monitor.scala 259:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_325 & ~_T_1384) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:260 assert (source_ok, \"'C' channel HintAck carries invalid source ID\" + extra)\n"); // @[Monitor.scala 260:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_325 & ~_T_1384) begin
          $fatal; // @[Monitor.scala 260:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_325 & ~_T_1391) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:261 assert (is_aligned, \"'C' channel HintAck address not aligned to size\" + extra)\n"); // @[Monitor.scala 261:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_325 & ~_T_1391) begin
          $fatal; // @[Monitor.scala 261:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_325 & ~_T_1617) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:262 assert (bundle.param === UInt(0), \"'C' channel HintAck carries invalid param\" + extra)\n"); // @[Monitor.scala 262:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_325 & ~_T_1617) begin
          $fatal; // @[Monitor.scala 262:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1692 & ~_T_1695) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:355 assert (a.bits.opcode === opcode, \"'A' channel opcode changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 355:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1692 & ~_T_1695) begin
          $fatal; // @[Monitor.scala 355:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1692 & ~_T_1699) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:356 assert (a.bits.param  === param,  \"'A' channel param changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 356:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1692 & ~_T_1699) begin
          $fatal; // @[Monitor.scala 356:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1692 & ~_T_1703) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:357 assert (a.bits.size   === size,   \"'A' channel size changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 357:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1692 & ~_T_1703) begin
          $fatal; // @[Monitor.scala 357:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1692 & ~_T_1707) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:358 assert (a.bits.source === source, \"'A' channel source changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 358:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1692 & ~_T_1707) begin
          $fatal; // @[Monitor.scala 358:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1692 & ~_T_1711) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:359 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); // @[Monitor.scala 359:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1692 & ~_T_1711) begin
          $fatal; // @[Monitor.scala 359:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1749 & ~_T_1752) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:425 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 425:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1749 & ~_T_1752) begin
          $fatal; // @[Monitor.scala 425:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1749 & ~_T_1756) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:426 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 426:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1749 & ~_T_1756) begin
          $fatal; // @[Monitor.scala 426:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1749 & ~_T_1760) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:427 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 427:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1749 & ~_T_1760) begin
          $fatal; // @[Monitor.scala 427:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1749 & ~_T_1764) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:428 assert (d.bits.source === source, \"'D' channel source changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 428:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1749 & ~_T_1764) begin
          $fatal; // @[Monitor.scala 428:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1749 & ~_T_1768) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:429 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); // @[Monitor.scala 429:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1749 & ~_T_1768) begin
          $fatal; // @[Monitor.scala 429:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1749 & ~_T_1772) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:430 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); // @[Monitor.scala 430:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1749 & ~_T_1772) begin
          $fatal; // @[Monitor.scala 430:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1809 & ~_T_1812) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel opcode changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:378 assert (b.bits.opcode === opcode, \"'B' channel opcode changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 378:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1809 & ~_T_1812) begin
          $fatal; // @[Monitor.scala 378:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1809 & ~_T_1816) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel param changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:379 assert (b.bits.param  === param,  \"'B' channel param changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 379:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1809 & ~_T_1816) begin
          $fatal; // @[Monitor.scala 379:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1809 & ~_T_1820) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel size changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:380 assert (b.bits.size   === size,   \"'B' channel size changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 380:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1809 & ~_T_1820) begin
          $fatal; // @[Monitor.scala 380:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1809 & ~_T_1824) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel source changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:381 assert (b.bits.source === source, \"'B' channel source changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 381:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1809 & ~_T_1824) begin
          $fatal; // @[Monitor.scala 381:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1809 & ~_T_1828) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel addresss changed with multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:382 assert (b.bits.address=== address,\"'B' channel addresss changed with multibeat operation\" + extra)\n"); // @[Monitor.scala 382:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1809 & ~_T_1828) begin
          $fatal; // @[Monitor.scala 382:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1864 & ~_T_1867) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel opcode changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:401 assert (c.bits.opcode === opcode, \"'C' channel opcode changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 401:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1864 & ~_T_1867) begin
          $fatal; // @[Monitor.scala 401:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1864 & ~_T_1871) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel param changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:402 assert (c.bits.param  === param,  \"'C' channel param changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 402:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1864 & ~_T_1871) begin
          $fatal; // @[Monitor.scala 402:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1864 & ~_T_1875) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel size changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:403 assert (c.bits.size   === size,   \"'C' channel size changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 403:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1864 & ~_T_1875) begin
          $fatal; // @[Monitor.scala 403:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1864 & ~_T_1879) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel source changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:404 assert (c.bits.source === source, \"'C' channel source changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 404:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1864 & ~_T_1879) begin
          $fatal; // @[Monitor.scala 404:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1864 & ~_T_1883) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel address changed with multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:405 assert (c.bits.address=== address,\"'C' channel address changed with multibeat operation\" + extra)\n"); // @[Monitor.scala 405:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1864 & ~_T_1883) begin
          $fatal; // @[Monitor.scala 405:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1935 & ~_T_1942) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:460 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); // @[Monitor.scala 460:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1935 & ~_T_1942) begin
          $fatal; // @[Monitor.scala 460:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1951 & ~_T_1957) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:467 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); // @[Monitor.scala 467:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1951 & ~_T_1957) begin
          $fatal; // @[Monitor.scala 467:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_1964) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:471 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); // @[Monitor.scala 471:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_1964) begin
          $fatal; // @[Monitor.scala 471:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2016 & ~_T_2022) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel re-used a sink ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:494 assert(!inflight(bundle.d.bits.sink), \"'D' channel re-used a sink ID\" + extra)\n"); // @[Monitor.scala 494:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2016 & ~_T_2022) begin
          $fatal; // @[Monitor.scala 494:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2026 & ~_T_2034) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel acknowledged for nothing inflight (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:500 assert((d_set | inflight)(bundle.e.bits.sink), \"'E' channel acknowledged for nothing inflight\" + extra)\n"); // @[Monitor.scala 500:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2026 & ~_T_2034) begin
          $fatal; // @[Monitor.scala 500:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    if (metaReset) begin
      TLMonitor_66_metaAssert <= 1'h0;
    end else begin
      TLMonitor_66_metaAssert <= TLMonitor_66_metaAssert | TLMonitor_66_or0;
    end
  end
endmodule
module Queue_108(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_param,
  input  [3:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_source,
  input  [31:0] io_enq_bits_address,
  input  [7:0]  io_enq_bits_mask,
  input  [63:0] io_enq_bits_data,
  input         io_enq_bits_corrupt,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_param,
  output [3:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_source,
  output [31:0] io_deq_bits_address,
  output [7:0]  io_deq_bits_mask,
  output [63:0] io_deq_bits_data,
  output        io_deq_bits_corrupt,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [2:0] _T_35_opcode [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_0;
  wire [2:0] _T_35_opcode__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_opcode__T_58_addr; // @[Decoupled.scala 214:24]
  wire [2:0] _T_35_opcode__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_opcode__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_opcode__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_opcode__T_50_en; // @[Decoupled.scala 214:24]
  reg [2:0] _T_35_param [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_1;
  wire [2:0] _T_35_param__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_param__T_58_addr; // @[Decoupled.scala 214:24]
  wire [2:0] _T_35_param__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_param__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_param__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_param__T_50_en; // @[Decoupled.scala 214:24]
  reg [3:0] _T_35_size [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_2;
  wire [3:0] _T_35_size__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_size__T_58_addr; // @[Decoupled.scala 214:24]
  wire [3:0] _T_35_size__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_size__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_size__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_size__T_50_en; // @[Decoupled.scala 214:24]
  reg [1:0] _T_35_source [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_3;
  wire [1:0] _T_35_source__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_source__T_58_addr; // @[Decoupled.scala 214:24]
  wire [1:0] _T_35_source__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_source__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_source__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_source__T_50_en; // @[Decoupled.scala 214:24]
  reg [31:0] _T_35_address [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_4;
  wire [31:0] _T_35_address__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_address__T_58_addr; // @[Decoupled.scala 214:24]
  wire [31:0] _T_35_address__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_address__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_address__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_address__T_50_en; // @[Decoupled.scala 214:24]
  reg [7:0] _T_35_mask [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_5;
  wire [7:0] _T_35_mask__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_mask__T_58_addr; // @[Decoupled.scala 214:24]
  wire [7:0] _T_35_mask__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_mask__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_mask__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_mask__T_50_en; // @[Decoupled.scala 214:24]
  reg [63:0] _T_35_data [0:1]; // @[Decoupled.scala 214:24]
  reg [63:0] _RAND_6;
  wire [63:0] _T_35_data__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_data__T_58_addr; // @[Decoupled.scala 214:24]
  wire [63:0] _T_35_data__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_data__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_data__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_data__T_50_en; // @[Decoupled.scala 214:24]
  reg  _T_35_corrupt [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_7;
  wire  _T_35_corrupt__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_corrupt__T_58_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_corrupt__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_corrupt__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_corrupt__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_corrupt__T_50_en; // @[Decoupled.scala 214:24]
  reg  value; // @[Counter.scala 26:33]
  reg [31:0] _RAND_8;
  reg  value_1; // @[Counter.scala 26:33]
  reg [31:0] _RAND_9;
  reg  _T_39; // @[Decoupled.scala 217:35]
  reg [31:0] _RAND_10;
  wire  _T_40; // @[Decoupled.scala 219:41]
  wire  _T_42; // @[Decoupled.scala 220:33]
  wire  _T_43; // @[Decoupled.scala 221:32]
  wire  _T_44; // @[Decoupled.scala 37:37]
  wire  _T_47; // @[Decoupled.scala 37:37]
  wire  _T_52; // @[Counter.scala 35:22]
  wire  _T_54; // @[Counter.scala 35:22]
  wire  _T_55; // @[Decoupled.scala 232:16]
  wire [29:0] Queue_108_covSum;
  assign _T_35_opcode__T_58_addr = value_1;
  assign _T_35_opcode__T_58_data = _T_35_opcode[_T_35_opcode__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_opcode__T_50_data = io_enq_bits_opcode;
  assign _T_35_opcode__T_50_addr = value;
  assign _T_35_opcode__T_50_mask = 1'h1;
  assign _T_35_opcode__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_param__T_58_addr = value_1;
  assign _T_35_param__T_58_data = _T_35_param[_T_35_param__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_param__T_50_data = io_enq_bits_param;
  assign _T_35_param__T_50_addr = value;
  assign _T_35_param__T_50_mask = 1'h1;
  assign _T_35_param__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_size__T_58_addr = value_1;
  assign _T_35_size__T_58_data = _T_35_size[_T_35_size__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_size__T_50_data = io_enq_bits_size;
  assign _T_35_size__T_50_addr = value;
  assign _T_35_size__T_50_mask = 1'h1;
  assign _T_35_size__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_source__T_58_addr = value_1;
  assign _T_35_source__T_58_data = _T_35_source[_T_35_source__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_source__T_50_data = io_enq_bits_source;
  assign _T_35_source__T_50_addr = value;
  assign _T_35_source__T_50_mask = 1'h1;
  assign _T_35_source__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_address__T_58_addr = value_1;
  assign _T_35_address__T_58_data = _T_35_address[_T_35_address__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_address__T_50_data = io_enq_bits_address;
  assign _T_35_address__T_50_addr = value;
  assign _T_35_address__T_50_mask = 1'h1;
  assign _T_35_address__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_mask__T_58_addr = value_1;
  assign _T_35_mask__T_58_data = _T_35_mask[_T_35_mask__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_mask__T_50_data = io_enq_bits_mask;
  assign _T_35_mask__T_50_addr = value;
  assign _T_35_mask__T_50_mask = 1'h1;
  assign _T_35_mask__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_data__T_58_addr = value_1;
  assign _T_35_data__T_58_data = _T_35_data[_T_35_data__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_data__T_50_data = io_enq_bits_data;
  assign _T_35_data__T_50_addr = value;
  assign _T_35_data__T_50_mask = 1'h1;
  assign _T_35_data__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_corrupt__T_58_addr = value_1;
  assign _T_35_corrupt__T_58_data = _T_35_corrupt[_T_35_corrupt__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_corrupt__T_50_data = io_enq_bits_corrupt;
  assign _T_35_corrupt__T_50_addr = value;
  assign _T_35_corrupt__T_50_mask = 1'h1;
  assign _T_35_corrupt__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_40 = value == value_1; // @[Decoupled.scala 219:41]
  assign _T_42 = _T_40 & ~_T_39; // @[Decoupled.scala 220:33]
  assign _T_43 = _T_40 & _T_39; // @[Decoupled.scala 221:32]
  assign _T_44 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37]
  assign _T_47 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 37:37]
  assign _T_52 = value + 1'h1; // @[Counter.scala 35:22]
  assign _T_54 = value_1 + 1'h1; // @[Counter.scala 35:22]
  assign _T_55 = _T_44 != _T_47; // @[Decoupled.scala 232:16]
  assign io_enq_ready = ~_T_43; // @[Decoupled.scala 237:16]
  assign io_deq_valid = ~_T_42; // @[Decoupled.scala 236:16]
  assign io_deq_bits_opcode = _T_35_opcode__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_param = _T_35_param__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_size = _T_35_size__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_source = _T_35_source__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_address = _T_35_address__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_mask = _T_35_mask__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_data = _T_35_data__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_corrupt = _T_35_corrupt__T_58_data; // @[Decoupled.scala 238:15]
  assign Queue_108_covSum = 30'h0;
  assign io_covSum = Queue_108_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_param[initvar] = _RAND_1[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_size[initvar] = _RAND_2[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_source[initvar] = _RAND_3[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_address[initvar] = _RAND_4[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_mask[initvar] = _RAND_5[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_data[initvar] = _RAND_6[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_corrupt[initvar] = _RAND_7[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_39 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_35_opcode__T_50_en & _T_35_opcode__T_50_mask) begin
      _T_35_opcode[_T_35_opcode__T_50_addr] <= _T_35_opcode__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_param__T_50_en & _T_35_param__T_50_mask) begin
      _T_35_param[_T_35_param__T_50_addr] <= _T_35_param__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_size__T_50_en & _T_35_size__T_50_mask) begin
      _T_35_size[_T_35_size__T_50_addr] <= _T_35_size__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_source__T_50_en & _T_35_source__T_50_mask) begin
      _T_35_source[_T_35_source__T_50_addr] <= _T_35_source__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_address__T_50_en & _T_35_address__T_50_mask) begin
      _T_35_address[_T_35_address__T_50_addr] <= _T_35_address__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_mask__T_50_en & _T_35_mask__T_50_mask) begin
      _T_35_mask[_T_35_mask__T_50_addr] <= _T_35_mask__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_data__T_50_en & _T_35_data__T_50_mask) begin
      _T_35_data[_T_35_data__T_50_addr] <= _T_35_data__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_corrupt__T_50_en & _T_35_corrupt__T_50_mask) begin
      _T_35_corrupt[_T_35_corrupt__T_50_addr] <= _T_35_corrupt__T_50_data; // @[Decoupled.scala 214:24]
    end
    if (metaReset) begin
      value <= 1'h0;
    end else if (reset) begin
      value <= 1'h0;
    end else if (_T_44) begin
      value <= _T_52;
    end
    if (metaReset) begin
      value_1 <= 1'h0;
    end else if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_47) begin
      value_1 <= _T_54;
    end
    if (metaReset) begin
      _T_39 <= 1'h0;
    end else if (reset) begin
      _T_39 <= 1'h0;
    end else if (_T_55) begin
      _T_39 <= _T_44;
    end
  end
endmodule
module Queue_109(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [1:0]  io_enq_bits_param,
  input  [3:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_source,
  input  [1:0]  io_enq_bits_sink,
  input         io_enq_bits_denied,
  input  [63:0] io_enq_bits_data,
  input         io_enq_bits_corrupt,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [1:0]  io_deq_bits_param,
  output [3:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_source,
  output [1:0]  io_deq_bits_sink,
  output        io_deq_bits_denied,
  output [63:0] io_deq_bits_data,
  output        io_deq_bits_corrupt,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [2:0] _T_35_opcode [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_0;
  wire [2:0] _T_35_opcode__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_opcode__T_58_addr; // @[Decoupled.scala 214:24]
  wire [2:0] _T_35_opcode__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_opcode__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_opcode__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_opcode__T_50_en; // @[Decoupled.scala 214:24]
  reg [1:0] _T_35_param [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_1;
  wire [1:0] _T_35_param__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_param__T_58_addr; // @[Decoupled.scala 214:24]
  wire [1:0] _T_35_param__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_param__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_param__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_param__T_50_en; // @[Decoupled.scala 214:24]
  reg [3:0] _T_35_size [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_2;
  wire [3:0] _T_35_size__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_size__T_58_addr; // @[Decoupled.scala 214:24]
  wire [3:0] _T_35_size__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_size__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_size__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_size__T_50_en; // @[Decoupled.scala 214:24]
  reg [1:0] _T_35_source [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_3;
  wire [1:0] _T_35_source__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_source__T_58_addr; // @[Decoupled.scala 214:24]
  wire [1:0] _T_35_source__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_source__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_source__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_source__T_50_en; // @[Decoupled.scala 214:24]
  reg [1:0] _T_35_sink [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_4;
  wire [1:0] _T_35_sink__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_sink__T_58_addr; // @[Decoupled.scala 214:24]
  wire [1:0] _T_35_sink__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_sink__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_sink__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_sink__T_50_en; // @[Decoupled.scala 214:24]
  reg  _T_35_denied [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_5;
  wire  _T_35_denied__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_denied__T_58_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_denied__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_denied__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_denied__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_denied__T_50_en; // @[Decoupled.scala 214:24]
  reg [63:0] _T_35_data [0:1]; // @[Decoupled.scala 214:24]
  reg [63:0] _RAND_6;
  wire [63:0] _T_35_data__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_data__T_58_addr; // @[Decoupled.scala 214:24]
  wire [63:0] _T_35_data__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_data__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_data__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_data__T_50_en; // @[Decoupled.scala 214:24]
  reg  _T_35_corrupt [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_7;
  wire  _T_35_corrupt__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_corrupt__T_58_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_corrupt__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_corrupt__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_corrupt__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_corrupt__T_50_en; // @[Decoupled.scala 214:24]
  reg  value; // @[Counter.scala 26:33]
  reg [31:0] _RAND_8;
  reg  value_1; // @[Counter.scala 26:33]
  reg [31:0] _RAND_9;
  reg  _T_39; // @[Decoupled.scala 217:35]
  reg [31:0] _RAND_10;
  wire  _T_40; // @[Decoupled.scala 219:41]
  wire  _T_42; // @[Decoupled.scala 220:33]
  wire  _T_43; // @[Decoupled.scala 221:32]
  wire  _T_44; // @[Decoupled.scala 37:37]
  wire  _T_47; // @[Decoupled.scala 37:37]
  wire  _T_52; // @[Counter.scala 35:22]
  wire  _T_54; // @[Counter.scala 35:22]
  wire  _T_55; // @[Decoupled.scala 232:16]
  wire [29:0] Queue_109_covSum;
  assign _T_35_opcode__T_58_addr = value_1;
  assign _T_35_opcode__T_58_data = _T_35_opcode[_T_35_opcode__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_opcode__T_50_data = io_enq_bits_opcode;
  assign _T_35_opcode__T_50_addr = value;
  assign _T_35_opcode__T_50_mask = 1'h1;
  assign _T_35_opcode__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_param__T_58_addr = value_1;
  assign _T_35_param__T_58_data = _T_35_param[_T_35_param__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_param__T_50_data = io_enq_bits_param;
  assign _T_35_param__T_50_addr = value;
  assign _T_35_param__T_50_mask = 1'h1;
  assign _T_35_param__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_size__T_58_addr = value_1;
  assign _T_35_size__T_58_data = _T_35_size[_T_35_size__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_size__T_50_data = io_enq_bits_size;
  assign _T_35_size__T_50_addr = value;
  assign _T_35_size__T_50_mask = 1'h1;
  assign _T_35_size__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_source__T_58_addr = value_1;
  assign _T_35_source__T_58_data = _T_35_source[_T_35_source__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_source__T_50_data = io_enq_bits_source;
  assign _T_35_source__T_50_addr = value;
  assign _T_35_source__T_50_mask = 1'h1;
  assign _T_35_source__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_sink__T_58_addr = value_1;
  assign _T_35_sink__T_58_data = _T_35_sink[_T_35_sink__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_sink__T_50_data = io_enq_bits_sink;
  assign _T_35_sink__T_50_addr = value;
  assign _T_35_sink__T_50_mask = 1'h1;
  assign _T_35_sink__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_denied__T_58_addr = value_1;
  assign _T_35_denied__T_58_data = _T_35_denied[_T_35_denied__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_denied__T_50_data = io_enq_bits_denied;
  assign _T_35_denied__T_50_addr = value;
  assign _T_35_denied__T_50_mask = 1'h1;
  assign _T_35_denied__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_data__T_58_addr = value_1;
  assign _T_35_data__T_58_data = _T_35_data[_T_35_data__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_data__T_50_data = io_enq_bits_data;
  assign _T_35_data__T_50_addr = value;
  assign _T_35_data__T_50_mask = 1'h1;
  assign _T_35_data__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_corrupt__T_58_addr = value_1;
  assign _T_35_corrupt__T_58_data = _T_35_corrupt[_T_35_corrupt__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_corrupt__T_50_data = io_enq_bits_corrupt;
  assign _T_35_corrupt__T_50_addr = value;
  assign _T_35_corrupt__T_50_mask = 1'h1;
  assign _T_35_corrupt__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_40 = value == value_1; // @[Decoupled.scala 219:41]
  assign _T_42 = _T_40 & ~_T_39; // @[Decoupled.scala 220:33]
  assign _T_43 = _T_40 & _T_39; // @[Decoupled.scala 221:32]
  assign _T_44 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37]
  assign _T_47 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 37:37]
  assign _T_52 = value + 1'h1; // @[Counter.scala 35:22]
  assign _T_54 = value_1 + 1'h1; // @[Counter.scala 35:22]
  assign _T_55 = _T_44 != _T_47; // @[Decoupled.scala 232:16]
  assign io_enq_ready = ~_T_43; // @[Decoupled.scala 237:16]
  assign io_deq_valid = ~_T_42; // @[Decoupled.scala 236:16]
  assign io_deq_bits_opcode = _T_35_opcode__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_param = _T_35_param__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_size = _T_35_size__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_source = _T_35_source__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_sink = _T_35_sink__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_denied = _T_35_denied__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_data = _T_35_data__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_corrupt = _T_35_corrupt__T_58_data; // @[Decoupled.scala 238:15]
  assign Queue_109_covSum = 30'h0;
  assign io_covSum = Queue_109_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_param[initvar] = _RAND_1[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_size[initvar] = _RAND_2[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_source[initvar] = _RAND_3[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_sink[initvar] = _RAND_4[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_denied[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_data[initvar] = _RAND_6[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_corrupt[initvar] = _RAND_7[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_39 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_35_opcode__T_50_en & _T_35_opcode__T_50_mask) begin
      _T_35_opcode[_T_35_opcode__T_50_addr] <= _T_35_opcode__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_param__T_50_en & _T_35_param__T_50_mask) begin
      _T_35_param[_T_35_param__T_50_addr] <= _T_35_param__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_size__T_50_en & _T_35_size__T_50_mask) begin
      _T_35_size[_T_35_size__T_50_addr] <= _T_35_size__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_source__T_50_en & _T_35_source__T_50_mask) begin
      _T_35_source[_T_35_source__T_50_addr] <= _T_35_source__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_sink__T_50_en & _T_35_sink__T_50_mask) begin
      _T_35_sink[_T_35_sink__T_50_addr] <= _T_35_sink__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_denied__T_50_en & _T_35_denied__T_50_mask) begin
      _T_35_denied[_T_35_denied__T_50_addr] <= _T_35_denied__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_data__T_50_en & _T_35_data__T_50_mask) begin
      _T_35_data[_T_35_data__T_50_addr] <= _T_35_data__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_corrupt__T_50_en & _T_35_corrupt__T_50_mask) begin
      _T_35_corrupt[_T_35_corrupt__T_50_addr] <= _T_35_corrupt__T_50_data; // @[Decoupled.scala 214:24]
    end
    if (metaReset) begin
      value <= 1'h0;
    end else if (reset) begin
      value <= 1'h0;
    end else if (_T_44) begin
      value <= _T_52;
    end
    if (metaReset) begin
      value_1 <= 1'h0;
    end else if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_47) begin
      value_1 <= _T_54;
    end
    if (metaReset) begin
      _T_39 <= 1'h0;
    end else if (reset) begin
      _T_39 <= 1'h0;
    end else if (_T_55) begin
      _T_39 <= _T_44;
    end
  end
endmodule
module Queue_110(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [1:0]  io_enq_bits_param,
  input  [3:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_source,
  input  [31:0] io_enq_bits_address,
  input  [7:0]  io_enq_bits_mask,
  input         io_enq_bits_corrupt,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [1:0]  io_deq_bits_param,
  output [3:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_source,
  output [31:0] io_deq_bits_address,
  output [7:0]  io_deq_bits_mask,
  output        io_deq_bits_corrupt,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [2:0] _T_35_opcode [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_0;
  wire [2:0] _T_35_opcode__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_opcode__T_58_addr; // @[Decoupled.scala 214:24]
  wire [2:0] _T_35_opcode__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_opcode__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_opcode__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_opcode__T_50_en; // @[Decoupled.scala 214:24]
  reg [1:0] _T_35_param [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_1;
  wire [1:0] _T_35_param__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_param__T_58_addr; // @[Decoupled.scala 214:24]
  wire [1:0] _T_35_param__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_param__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_param__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_param__T_50_en; // @[Decoupled.scala 214:24]
  reg [3:0] _T_35_size [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_2;
  wire [3:0] _T_35_size__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_size__T_58_addr; // @[Decoupled.scala 214:24]
  wire [3:0] _T_35_size__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_size__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_size__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_size__T_50_en; // @[Decoupled.scala 214:24]
  reg [1:0] _T_35_source [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_3;
  wire [1:0] _T_35_source__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_source__T_58_addr; // @[Decoupled.scala 214:24]
  wire [1:0] _T_35_source__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_source__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_source__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_source__T_50_en; // @[Decoupled.scala 214:24]
  reg [31:0] _T_35_address [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_4;
  wire [31:0] _T_35_address__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_address__T_58_addr; // @[Decoupled.scala 214:24]
  wire [31:0] _T_35_address__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_address__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_address__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_address__T_50_en; // @[Decoupled.scala 214:24]
  reg [7:0] _T_35_mask [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_5;
  wire [7:0] _T_35_mask__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_mask__T_58_addr; // @[Decoupled.scala 214:24]
  wire [7:0] _T_35_mask__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_mask__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_mask__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_mask__T_50_en; // @[Decoupled.scala 214:24]
  reg  _T_35_corrupt [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_6;
  wire  _T_35_corrupt__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_corrupt__T_58_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_corrupt__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_corrupt__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_corrupt__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_corrupt__T_50_en; // @[Decoupled.scala 214:24]
  reg  value; // @[Counter.scala 26:33]
  reg [31:0] _RAND_7;
  reg  value_1; // @[Counter.scala 26:33]
  reg [31:0] _RAND_8;
  reg  _T_39; // @[Decoupled.scala 217:35]
  reg [31:0] _RAND_9;
  wire  _T_40; // @[Decoupled.scala 219:41]
  wire  _T_42; // @[Decoupled.scala 220:33]
  wire  _T_43; // @[Decoupled.scala 221:32]
  wire  _T_44; // @[Decoupled.scala 37:37]
  wire  _T_47; // @[Decoupled.scala 37:37]
  wire  _T_52; // @[Counter.scala 35:22]
  wire  _T_54; // @[Counter.scala 35:22]
  wire  _T_55; // @[Decoupled.scala 232:16]
  wire [29:0] Queue_110_covSum;
  assign _T_35_opcode__T_58_addr = value_1;
  assign _T_35_opcode__T_58_data = _T_35_opcode[_T_35_opcode__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_opcode__T_50_data = io_enq_bits_opcode;
  assign _T_35_opcode__T_50_addr = value;
  assign _T_35_opcode__T_50_mask = 1'h1;
  assign _T_35_opcode__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_param__T_58_addr = value_1;
  assign _T_35_param__T_58_data = _T_35_param[_T_35_param__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_param__T_50_data = io_enq_bits_param;
  assign _T_35_param__T_50_addr = value;
  assign _T_35_param__T_50_mask = 1'h1;
  assign _T_35_param__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_size__T_58_addr = value_1;
  assign _T_35_size__T_58_data = _T_35_size[_T_35_size__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_size__T_50_data = io_enq_bits_size;
  assign _T_35_size__T_50_addr = value;
  assign _T_35_size__T_50_mask = 1'h1;
  assign _T_35_size__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_source__T_58_addr = value_1;
  assign _T_35_source__T_58_data = _T_35_source[_T_35_source__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_source__T_50_data = io_enq_bits_source;
  assign _T_35_source__T_50_addr = value;
  assign _T_35_source__T_50_mask = 1'h1;
  assign _T_35_source__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_address__T_58_addr = value_1;
  assign _T_35_address__T_58_data = _T_35_address[_T_35_address__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_address__T_50_data = io_enq_bits_address;
  assign _T_35_address__T_50_addr = value;
  assign _T_35_address__T_50_mask = 1'h1;
  assign _T_35_address__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_mask__T_58_addr = value_1;
  assign _T_35_mask__T_58_data = _T_35_mask[_T_35_mask__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_mask__T_50_data = io_enq_bits_mask;
  assign _T_35_mask__T_50_addr = value;
  assign _T_35_mask__T_50_mask = 1'h1;
  assign _T_35_mask__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_corrupt__T_58_addr = value_1;
  assign _T_35_corrupt__T_58_data = _T_35_corrupt[_T_35_corrupt__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_corrupt__T_50_data = io_enq_bits_corrupt;
  assign _T_35_corrupt__T_50_addr = value;
  assign _T_35_corrupt__T_50_mask = 1'h1;
  assign _T_35_corrupt__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_40 = value == value_1; // @[Decoupled.scala 219:41]
  assign _T_42 = _T_40 & ~_T_39; // @[Decoupled.scala 220:33]
  assign _T_43 = _T_40 & _T_39; // @[Decoupled.scala 221:32]
  assign _T_44 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37]
  assign _T_47 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 37:37]
  assign _T_52 = value + 1'h1; // @[Counter.scala 35:22]
  assign _T_54 = value_1 + 1'h1; // @[Counter.scala 35:22]
  assign _T_55 = _T_44 != _T_47; // @[Decoupled.scala 232:16]
  assign io_enq_ready = ~_T_43; // @[Decoupled.scala 237:16]
  assign io_deq_valid = ~_T_42; // @[Decoupled.scala 236:16]
  assign io_deq_bits_opcode = _T_35_opcode__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_param = _T_35_param__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_size = _T_35_size__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_source = _T_35_source__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_address = _T_35_address__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_mask = _T_35_mask__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_corrupt = _T_35_corrupt__T_58_data; // @[Decoupled.scala 238:15]
  assign Queue_110_covSum = 30'h0;
  assign io_covSum = Queue_110_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_param[initvar] = _RAND_1[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_size[initvar] = _RAND_2[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_source[initvar] = _RAND_3[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_address[initvar] = _RAND_4[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_mask[initvar] = _RAND_5[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_corrupt[initvar] = _RAND_6[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value_1 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_39 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_35_opcode__T_50_en & _T_35_opcode__T_50_mask) begin
      _T_35_opcode[_T_35_opcode__T_50_addr] <= _T_35_opcode__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_param__T_50_en & _T_35_param__T_50_mask) begin
      _T_35_param[_T_35_param__T_50_addr] <= _T_35_param__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_size__T_50_en & _T_35_size__T_50_mask) begin
      _T_35_size[_T_35_size__T_50_addr] <= _T_35_size__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_source__T_50_en & _T_35_source__T_50_mask) begin
      _T_35_source[_T_35_source__T_50_addr] <= _T_35_source__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_address__T_50_en & _T_35_address__T_50_mask) begin
      _T_35_address[_T_35_address__T_50_addr] <= _T_35_address__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_mask__T_50_en & _T_35_mask__T_50_mask) begin
      _T_35_mask[_T_35_mask__T_50_addr] <= _T_35_mask__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_corrupt__T_50_en & _T_35_corrupt__T_50_mask) begin
      _T_35_corrupt[_T_35_corrupt__T_50_addr] <= _T_35_corrupt__T_50_data; // @[Decoupled.scala 214:24]
    end
    if (metaReset) begin
      value <= 1'h0;
    end else if (reset) begin
      value <= 1'h0;
    end else if (_T_44) begin
      value <= _T_52;
    end
    if (metaReset) begin
      value_1 <= 1'h0;
    end else if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_47) begin
      value_1 <= _T_54;
    end
    if (metaReset) begin
      _T_39 <= 1'h0;
    end else if (reset) begin
      _T_39 <= 1'h0;
    end else if (_T_55) begin
      _T_39 <= _T_44;
    end
  end
endmodule
module Queue_111(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_param,
  input  [3:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_source,
  input  [31:0] io_enq_bits_address,
  input  [63:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_param,
  output [3:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_source,
  output [31:0] io_deq_bits_address,
  output [63:0] io_deq_bits_data,
  output        io_deq_bits_corrupt,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [2:0] _T_35_opcode [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_0;
  wire [2:0] _T_35_opcode__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_opcode__T_58_addr; // @[Decoupled.scala 214:24]
  wire [2:0] _T_35_opcode__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_opcode__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_opcode__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_opcode__T_50_en; // @[Decoupled.scala 214:24]
  reg [2:0] _T_35_param [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_1;
  wire [2:0] _T_35_param__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_param__T_58_addr; // @[Decoupled.scala 214:24]
  wire [2:0] _T_35_param__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_param__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_param__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_param__T_50_en; // @[Decoupled.scala 214:24]
  reg [3:0] _T_35_size [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_2;
  wire [3:0] _T_35_size__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_size__T_58_addr; // @[Decoupled.scala 214:24]
  wire [3:0] _T_35_size__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_size__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_size__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_size__T_50_en; // @[Decoupled.scala 214:24]
  reg [1:0] _T_35_source [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_3;
  wire [1:0] _T_35_source__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_source__T_58_addr; // @[Decoupled.scala 214:24]
  wire [1:0] _T_35_source__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_source__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_source__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_source__T_50_en; // @[Decoupled.scala 214:24]
  reg [31:0] _T_35_address [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_4;
  wire [31:0] _T_35_address__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_address__T_58_addr; // @[Decoupled.scala 214:24]
  wire [31:0] _T_35_address__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_address__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_address__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_address__T_50_en; // @[Decoupled.scala 214:24]
  reg [63:0] _T_35_data [0:1]; // @[Decoupled.scala 214:24]
  reg [63:0] _RAND_5;
  wire [63:0] _T_35_data__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_data__T_58_addr; // @[Decoupled.scala 214:24]
  wire [63:0] _T_35_data__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_data__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_data__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_data__T_50_en; // @[Decoupled.scala 214:24]
  reg  _T_35_corrupt [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_6;
  wire  _T_35_corrupt__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_corrupt__T_58_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_corrupt__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_corrupt__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_corrupt__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_corrupt__T_50_en; // @[Decoupled.scala 214:24]
  reg  value; // @[Counter.scala 26:33]
  reg [31:0] _RAND_7;
  reg  value_1; // @[Counter.scala 26:33]
  reg [31:0] _RAND_8;
  reg  _T_39; // @[Decoupled.scala 217:35]
  reg [31:0] _RAND_9;
  wire  _T_40; // @[Decoupled.scala 219:41]
  wire  _T_42; // @[Decoupled.scala 220:33]
  wire  _T_43; // @[Decoupled.scala 221:32]
  wire  _T_44; // @[Decoupled.scala 37:37]
  wire  _T_47; // @[Decoupled.scala 37:37]
  wire  _T_52; // @[Counter.scala 35:22]
  wire  _T_54; // @[Counter.scala 35:22]
  wire  _T_55; // @[Decoupled.scala 232:16]
  wire [29:0] Queue_111_covSum;
  assign _T_35_opcode__T_58_addr = value_1;
  assign _T_35_opcode__T_58_data = _T_35_opcode[_T_35_opcode__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_opcode__T_50_data = io_enq_bits_opcode;
  assign _T_35_opcode__T_50_addr = value;
  assign _T_35_opcode__T_50_mask = 1'h1;
  assign _T_35_opcode__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_param__T_58_addr = value_1;
  assign _T_35_param__T_58_data = _T_35_param[_T_35_param__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_param__T_50_data = io_enq_bits_param;
  assign _T_35_param__T_50_addr = value;
  assign _T_35_param__T_50_mask = 1'h1;
  assign _T_35_param__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_size__T_58_addr = value_1;
  assign _T_35_size__T_58_data = _T_35_size[_T_35_size__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_size__T_50_data = io_enq_bits_size;
  assign _T_35_size__T_50_addr = value;
  assign _T_35_size__T_50_mask = 1'h1;
  assign _T_35_size__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_source__T_58_addr = value_1;
  assign _T_35_source__T_58_data = _T_35_source[_T_35_source__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_source__T_50_data = io_enq_bits_source;
  assign _T_35_source__T_50_addr = value;
  assign _T_35_source__T_50_mask = 1'h1;
  assign _T_35_source__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_address__T_58_addr = value_1;
  assign _T_35_address__T_58_data = _T_35_address[_T_35_address__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_address__T_50_data = io_enq_bits_address;
  assign _T_35_address__T_50_addr = value;
  assign _T_35_address__T_50_mask = 1'h1;
  assign _T_35_address__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_data__T_58_addr = value_1;
  assign _T_35_data__T_58_data = _T_35_data[_T_35_data__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_data__T_50_data = io_enq_bits_data;
  assign _T_35_data__T_50_addr = value;
  assign _T_35_data__T_50_mask = 1'h1;
  assign _T_35_data__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_35_corrupt__T_58_addr = value_1;
  assign _T_35_corrupt__T_58_data = _T_35_corrupt[_T_35_corrupt__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_corrupt__T_50_data = 1'h0;
  assign _T_35_corrupt__T_50_addr = value;
  assign _T_35_corrupt__T_50_mask = 1'h1;
  assign _T_35_corrupt__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_40 = value == value_1; // @[Decoupled.scala 219:41]
  assign _T_42 = _T_40 & ~_T_39; // @[Decoupled.scala 220:33]
  assign _T_43 = _T_40 & _T_39; // @[Decoupled.scala 221:32]
  assign _T_44 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37]
  assign _T_47 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 37:37]
  assign _T_52 = value + 1'h1; // @[Counter.scala 35:22]
  assign _T_54 = value_1 + 1'h1; // @[Counter.scala 35:22]
  assign _T_55 = _T_44 != _T_47; // @[Decoupled.scala 232:16]
  assign io_enq_ready = ~_T_43; // @[Decoupled.scala 237:16]
  assign io_deq_valid = ~_T_42; // @[Decoupled.scala 236:16]
  assign io_deq_bits_opcode = _T_35_opcode__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_param = _T_35_param__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_size = _T_35_size__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_source = _T_35_source__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_address = _T_35_address__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_data = _T_35_data__T_58_data; // @[Decoupled.scala 238:15]
  assign io_deq_bits_corrupt = _T_35_corrupt__T_58_data; // @[Decoupled.scala 238:15]
  assign Queue_111_covSum = 30'h0;
  assign io_covSum = Queue_111_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_param[initvar] = _RAND_1[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_size[initvar] = _RAND_2[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_source[initvar] = _RAND_3[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_address[initvar] = _RAND_4[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_data[initvar] = _RAND_5[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_corrupt[initvar] = _RAND_6[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value_1 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_39 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_35_opcode__T_50_en & _T_35_opcode__T_50_mask) begin
      _T_35_opcode[_T_35_opcode__T_50_addr] <= _T_35_opcode__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_param__T_50_en & _T_35_param__T_50_mask) begin
      _T_35_param[_T_35_param__T_50_addr] <= _T_35_param__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_size__T_50_en & _T_35_size__T_50_mask) begin
      _T_35_size[_T_35_size__T_50_addr] <= _T_35_size__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_source__T_50_en & _T_35_source__T_50_mask) begin
      _T_35_source[_T_35_source__T_50_addr] <= _T_35_source__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_address__T_50_en & _T_35_address__T_50_mask) begin
      _T_35_address[_T_35_address__T_50_addr] <= _T_35_address__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_data__T_50_en & _T_35_data__T_50_mask) begin
      _T_35_data[_T_35_data__T_50_addr] <= _T_35_data__T_50_data; // @[Decoupled.scala 214:24]
    end
    if(_T_35_corrupt__T_50_en & _T_35_corrupt__T_50_mask) begin
      _T_35_corrupt[_T_35_corrupt__T_50_addr] <= _T_35_corrupt__T_50_data; // @[Decoupled.scala 214:24]
    end
    if (metaReset) begin
      value <= 1'h0;
    end else if (reset) begin
      value <= 1'h0;
    end else if (_T_44) begin
      value <= _T_52;
    end
    if (metaReset) begin
      value_1 <= 1'h0;
    end else if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_47) begin
      value_1 <= _T_54;
    end
    if (metaReset) begin
      _T_39 <= 1'h0;
    end else if (reset) begin
      _T_39 <= 1'h0;
    end else if (_T_55) begin
      _T_39 <= _T_44;
    end
  end
endmodule
module Queue_112(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [1:0]  io_enq_bits_sink,
  input         io_deq_ready,
  output        io_deq_valid,
  output [1:0]  io_deq_bits_sink,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [1:0] _T_35_sink [0:1]; // @[Decoupled.scala 214:24]
  reg [31:0] _RAND_0;
  wire [1:0] _T_35_sink__T_58_data; // @[Decoupled.scala 214:24]
  wire  _T_35_sink__T_58_addr; // @[Decoupled.scala 214:24]
  wire [1:0] _T_35_sink__T_50_data; // @[Decoupled.scala 214:24]
  wire  _T_35_sink__T_50_addr; // @[Decoupled.scala 214:24]
  wire  _T_35_sink__T_50_mask; // @[Decoupled.scala 214:24]
  wire  _T_35_sink__T_50_en; // @[Decoupled.scala 214:24]
  reg  value; // @[Counter.scala 26:33]
  reg [31:0] _RAND_1;
  reg  value_1; // @[Counter.scala 26:33]
  reg [31:0] _RAND_2;
  reg  _T_39; // @[Decoupled.scala 217:35]
  reg [31:0] _RAND_3;
  wire  _T_40; // @[Decoupled.scala 219:41]
  wire  _T_42; // @[Decoupled.scala 220:33]
  wire  _T_43; // @[Decoupled.scala 221:32]
  wire  _T_44; // @[Decoupled.scala 37:37]
  wire  _T_47; // @[Decoupled.scala 37:37]
  wire  _T_52; // @[Counter.scala 35:22]
  wire  _T_54; // @[Counter.scala 35:22]
  wire  _T_55; // @[Decoupled.scala 232:16]
  wire [29:0] Queue_112_covSum;
  assign _T_35_sink__T_58_addr = value_1;
  assign _T_35_sink__T_58_data = _T_35_sink[_T_35_sink__T_58_addr]; // @[Decoupled.scala 214:24]
  assign _T_35_sink__T_50_data = io_enq_bits_sink;
  assign _T_35_sink__T_50_addr = value;
  assign _T_35_sink__T_50_mask = 1'h1;
  assign _T_35_sink__T_50_en = io_enq_ready & io_enq_valid;
  assign _T_40 = value == value_1; // @[Decoupled.scala 219:41]
  assign _T_42 = _T_40 & ~_T_39; // @[Decoupled.scala 220:33]
  assign _T_43 = _T_40 & _T_39; // @[Decoupled.scala 221:32]
  assign _T_44 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37]
  assign _T_47 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 37:37]
  assign _T_52 = value + 1'h1; // @[Counter.scala 35:22]
  assign _T_54 = value_1 + 1'h1; // @[Counter.scala 35:22]
  assign _T_55 = _T_44 != _T_47; // @[Decoupled.scala 232:16]
  assign io_enq_ready = ~_T_43; // @[Decoupled.scala 237:16]
  assign io_deq_valid = ~_T_42; // @[Decoupled.scala 236:16]
  assign io_deq_bits_sink = _T_35_sink__T_58_data; // @[Decoupled.scala 238:15]
  assign Queue_112_covSum = 30'h0;
  assign io_covSum = Queue_112_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_35_sink[initvar] = _RAND_0[1:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_39 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_35_sink__T_50_en & _T_35_sink__T_50_mask) begin
      _T_35_sink[_T_35_sink__T_50_addr] <= _T_35_sink__T_50_data; // @[Decoupled.scala 214:24]
    end
    if (metaReset) begin
      value <= 1'h0;
    end else if (reset) begin
      value <= 1'h0;
    end else if (_T_44) begin
      value <= _T_52;
    end
    if (metaReset) begin
      value_1 <= 1'h0;
    end else if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_47) begin
      value_1 <= _T_54;
    end
    if (metaReset) begin
      _T_39 <= 1'h0;
    end else if (reset) begin
      _T_39 <= 1'h0;
    end else if (_T_55) begin
      _T_39 <= _T_44;
    end
  end
endmodule
module SynchronizerShiftReg_w1_d3(
  input         clock,
  input         io_d,
  output        io_q,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg  sync_0; // @[ShiftReg.scala 114:16]
  reg [31:0] _RAND_0;
  reg  sync_1; // @[ShiftReg.scala 114:16]
  reg [31:0] _RAND_1;
  reg  sync_2; // @[ShiftReg.scala 114:16]
  reg [31:0] _RAND_2;
  wire [29:0] SynchronizerShiftReg_w1_d3_covSum;
  assign io_q = sync_0; // @[ShiftReg.scala 123:8]
  assign SynchronizerShiftReg_w1_d3_covSum = 30'h0;
  assign io_covSum = SynchronizerShiftReg_w1_d3_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sync_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sync_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  sync_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      sync_0 <= 1'h0;
    end else begin
      sync_0 <= sync_1;
    end
    if (metaReset) begin
      sync_1 <= 1'h0;
    end else begin
      sync_1 <= sync_2;
    end
    if (metaReset) begin
      sync_2 <= 1'h0;
    end else begin
      sync_2 <= io_d;
    end
  end
endmodule
module FPUDecoder(
  input  [31:0] io_inst,
  output        io_sigs_wen,
  output        io_sigs_ren1,
  output        io_sigs_ren2,
  output        io_sigs_ren3,
  output        io_sigs_swap12,
  output        io_sigs_swap23,
  output        io_sigs_singleIn,
  output        io_sigs_singleOut,
  output        io_sigs_fromint,
  output        io_sigs_toint,
  output        io_sigs_fastpipe,
  output        io_sigs_fma,
  output        io_sigs_div,
  output        io_sigs_sqrt,
  output        io_sigs_wflags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [31:0] _T_6; // @[Decode.scala 14:65]
  wire [31:0] _T_8; // @[Decode.scala 14:65]
  wire  _T_9; // @[Decode.scala 14:121]
  wire [31:0] _T_10; // @[Decode.scala 14:65]
  wire  _T_11; // @[Decode.scala 14:121]
  wire [31:0] _T_12; // @[Decode.scala 14:65]
  wire  _T_13; // @[Decode.scala 14:121]
  wire  _T_15; // @[Decode.scala 15:30]
  wire [31:0] _T_16; // @[Decode.scala 14:65]
  wire  _T_17; // @[Decode.scala 14:121]
  wire [31:0] _T_18; // @[Decode.scala 14:65]
  wire  _T_19; // @[Decode.scala 14:121]
  wire [31:0] _T_20; // @[Decode.scala 14:65]
  wire  decoder_4; // @[Decode.scala 14:121]
  wire  _T_23; // @[Decode.scala 15:30]
  wire [31:0] _T_24; // @[Decode.scala 14:65]
  wire  _T_25; // @[Decode.scala 14:121]
  wire [31:0] _T_26; // @[Decode.scala 14:65]
  wire  _T_27; // @[Decode.scala 14:121]
  wire  _T_29; // @[Decode.scala 15:30]
  wire [31:0] _T_30; // @[Decode.scala 14:65]
  wire [31:0] _T_32; // @[Decode.scala 14:65]
  wire  _T_33; // @[Decode.scala 14:121]
  wire [31:0] _T_34; // @[Decode.scala 14:65]
  wire  _T_35; // @[Decode.scala 14:121]
  wire [31:0] _T_36; // @[Decode.scala 14:65]
  wire  _T_37; // @[Decode.scala 14:121]
  wire [31:0] _T_38; // @[Decode.scala 14:65]
  wire  _T_39; // @[Decode.scala 14:121]
  wire [31:0] _T_40; // @[Decode.scala 14:65]
  wire  _T_41; // @[Decode.scala 14:121]
  wire [31:0] _T_42; // @[Decode.scala 14:65]
  wire  _T_43; // @[Decode.scala 14:121]
  wire [31:0] _T_44; // @[Decode.scala 14:65]
  wire  _T_45; // @[Decode.scala 14:121]
  wire  _T_47; // @[Decode.scala 15:30]
  wire  _T_48; // @[Decode.scala 15:30]
  wire  _T_49; // @[Decode.scala 15:30]
  wire  _T_50; // @[Decode.scala 15:30]
  wire  _T_51; // @[Decode.scala 15:30]
  wire [31:0] _T_52; // @[Decode.scala 14:65]
  wire  _T_53; // @[Decode.scala 14:121]
  wire [31:0] _T_54; // @[Decode.scala 14:65]
  wire  _T_55; // @[Decode.scala 14:121]
  wire  _T_57; // @[Decode.scala 14:121]
  wire [31:0] _T_58; // @[Decode.scala 14:65]
  wire  _T_59; // @[Decode.scala 14:121]
  wire [31:0] _T_60; // @[Decode.scala 14:65]
  wire  _T_61; // @[Decode.scala 14:121]
  wire  _T_63; // @[Decode.scala 15:30]
  wire  _T_64; // @[Decode.scala 15:30]
  wire  _T_65; // @[Decode.scala 15:30]
  wire [31:0] _T_66; // @[Decode.scala 14:65]
  wire  _T_69; // @[Decode.scala 14:121]
  wire [31:0] _T_71; // @[Decode.scala 14:65]
  wire  _T_72; // @[Decode.scala 14:121]
  wire [31:0] _T_73; // @[Decode.scala 14:65]
  wire  _T_74; // @[Decode.scala 14:121]
  wire [31:0] _T_76; // @[Decode.scala 14:65]
  wire  _T_77; // @[Decode.scala 14:121]
  wire [31:0] _T_78; // @[Decode.scala 14:65]
  wire  _T_79; // @[Decode.scala 14:121]
  wire  _T_81; // @[Decode.scala 15:30]
  wire [31:0] _T_82; // @[Decode.scala 14:65]
  wire [31:0] _T_86; // @[Decode.scala 14:65]
  wire  _T_87; // @[Decode.scala 14:121]
  wire [31:0] _T_88; // @[Decode.scala 14:65]
  wire  _T_89; // @[Decode.scala 14:121]
  wire [31:0] _T_90; // @[Decode.scala 14:65]
  wire  _T_91; // @[Decode.scala 14:121]
  wire  _T_93; // @[Decode.scala 15:30]
  wire  _T_94; // @[Decode.scala 15:30]
  wire [29:0] FPUDecoder_covSum;
  assign _T_6 = io_inst & 32'h40; // @[Decode.scala 14:65]
  assign _T_8 = io_inst & 32'h80000020; // @[Decode.scala 14:65]
  assign _T_9 = _T_8 == 32'h0; // @[Decode.scala 14:121]
  assign _T_10 = io_inst & 32'h30; // @[Decode.scala 14:65]
  assign _T_11 = _T_10 == 32'h0; // @[Decode.scala 14:121]
  assign _T_12 = io_inst & 32'h10000020; // @[Decode.scala 14:65]
  assign _T_13 = _T_12 == 32'h10000000; // @[Decode.scala 14:121]
  assign _T_15 = _T_9 | _T_11; // @[Decode.scala 15:30]
  assign _T_16 = io_inst & 32'h80000004; // @[Decode.scala 14:65]
  assign _T_17 = _T_16 == 32'h0; // @[Decode.scala 14:121]
  assign _T_18 = io_inst & 32'h10000004; // @[Decode.scala 14:65]
  assign _T_19 = _T_18 == 32'h0; // @[Decode.scala 14:121]
  assign _T_20 = io_inst & 32'h50; // @[Decode.scala 14:65]
  assign decoder_4 = _T_20 == 32'h40; // @[Decode.scala 14:121]
  assign _T_23 = _T_17 | _T_19; // @[Decode.scala 15:30]
  assign _T_24 = io_inst & 32'h40000004; // @[Decode.scala 14:65]
  assign _T_25 = _T_24 == 32'h0; // @[Decode.scala 14:121]
  assign _T_26 = io_inst & 32'h20; // @[Decode.scala 14:65]
  assign _T_27 = _T_26 == 32'h20; // @[Decode.scala 14:121]
  assign _T_29 = _T_25 | _T_27; // @[Decode.scala 15:30]
  assign _T_30 = io_inst & 32'h30000010; // @[Decode.scala 14:65]
  assign _T_32 = io_inst & 32'h82100020; // @[Decode.scala 14:65]
  assign _T_33 = _T_32 == 32'h0; // @[Decode.scala 14:121]
  assign _T_34 = io_inst & 32'h42000020; // @[Decode.scala 14:65]
  assign _T_35 = _T_34 == 32'h0; // @[Decode.scala 14:121]
  assign _T_36 = io_inst & 32'h2000030; // @[Decode.scala 14:65]
  assign _T_37 = _T_36 == 32'h0; // @[Decode.scala 14:121]
  assign _T_38 = io_inst & 32'h2103000; // @[Decode.scala 14:65]
  assign _T_39 = _T_38 == 32'h1000; // @[Decode.scala 14:121]
  assign _T_40 = io_inst & 32'h12002000; // @[Decode.scala 14:65]
  assign _T_41 = _T_40 == 32'h10000000; // @[Decode.scala 14:121]
  assign _T_42 = io_inst & 32'hd0100010; // @[Decode.scala 14:65]
  assign _T_43 = _T_42 == 32'h40000010; // @[Decode.scala 14:121]
  assign _T_44 = io_inst & 32'ha2000020; // @[Decode.scala 14:65]
  assign _T_45 = _T_44 == 32'h80000000; // @[Decode.scala 14:121]
  assign _T_47 = _T_33 | _T_35; // @[Decode.scala 15:30]
  assign _T_48 = _T_47 | _T_37; // @[Decode.scala 15:30]
  assign _T_49 = _T_48 | _T_39; // @[Decode.scala 15:30]
  assign _T_50 = _T_49 | _T_41; // @[Decode.scala 15:30]
  assign _T_51 = _T_50 | _T_43; // @[Decode.scala 15:30]
  assign _T_52 = io_inst & 32'h42001000; // @[Decode.scala 14:65]
  assign _T_53 = _T_52 == 32'h0; // @[Decode.scala 14:121]
  assign _T_54 = io_inst & 32'h22000004; // @[Decode.scala 14:65]
  assign _T_55 = _T_54 == 32'h0; // @[Decode.scala 14:121]
  assign _T_57 = _T_40 == 32'h0; // @[Decode.scala 14:121]
  assign _T_58 = io_inst & 32'h1040; // @[Decode.scala 14:65]
  assign _T_59 = _T_58 == 32'h0; // @[Decode.scala 14:121]
  assign _T_60 = io_inst & 32'h2000050; // @[Decode.scala 14:65]
  assign _T_61 = _T_60 == 32'h40; // @[Decode.scala 14:121]
  assign _T_63 = _T_53 | _T_55; // @[Decode.scala 15:30]
  assign _T_64 = _T_63 | _T_57; // @[Decode.scala 15:30]
  assign _T_65 = _T_64 | _T_59; // @[Decode.scala 15:30]
  assign _T_66 = io_inst & 32'h90000010; // @[Decode.scala 14:65]
  assign _T_69 = _T_66 == 32'h80000010; // @[Decode.scala 14:121]
  assign _T_71 = io_inst & 32'ha0000010; // @[Decode.scala 14:65]
  assign _T_72 = _T_71 == 32'h20000010; // @[Decode.scala 14:121]
  assign _T_73 = io_inst & 32'hd0000010; // @[Decode.scala 14:65]
  assign _T_74 = _T_73 == 32'h40000010; // @[Decode.scala 14:121]
  assign _T_76 = io_inst & 32'h70000004; // @[Decode.scala 14:65]
  assign _T_77 = _T_76 == 32'h0; // @[Decode.scala 14:121]
  assign _T_78 = io_inst & 32'h68000004; // @[Decode.scala 14:65]
  assign _T_79 = _T_78 == 32'h0; // @[Decode.scala 14:121]
  assign _T_81 = _T_77 | _T_79; // @[Decode.scala 15:30]
  assign _T_82 = io_inst & 32'h58000010; // @[Decode.scala 14:65]
  assign _T_86 = io_inst & 32'h20000004; // @[Decode.scala 14:65]
  assign _T_87 = _T_86 == 32'h0; // @[Decode.scala 14:121]
  assign _T_88 = io_inst & 32'h8002000; // @[Decode.scala 14:65]
  assign _T_89 = _T_88 == 32'h8000000; // @[Decode.scala 14:121]
  assign _T_90 = io_inst & 32'hc0000004; // @[Decode.scala 14:65]
  assign _T_91 = _T_90 == 32'h80000000; // @[Decode.scala 14:121]
  assign _T_93 = _T_87 | decoder_4; // @[Decode.scala 15:30]
  assign _T_94 = _T_93 | _T_89; // @[Decode.scala 15:30]
  assign io_sigs_wen = _T_15 | _T_13; // @[FPU.scala 133:40]
  assign io_sigs_ren1 = _T_23 | decoder_4; // @[FPU.scala 133:40]
  assign io_sigs_ren2 = _T_29 | decoder_4; // @[FPU.scala 133:40]
  assign io_sigs_ren3 = _T_20 == 32'h40; // @[FPU.scala 133:40]
  assign io_sigs_swap12 = _T_6 == 32'h0; // @[FPU.scala 133:40]
  assign io_sigs_swap23 = _T_30 == 32'h10; // @[FPU.scala 133:40]
  assign io_sigs_singleIn = _T_51 | _T_45; // @[FPU.scala 133:40]
  assign io_sigs_singleOut = _T_65 | _T_61; // @[FPU.scala 133:40]
  assign io_sigs_fromint = _T_66 == 32'h90000010; // @[FPU.scala 133:40]
  assign io_sigs_toint = _T_27 | _T_69; // @[FPU.scala 133:40]
  assign io_sigs_fastpipe = _T_72 | _T_74; // @[FPU.scala 133:40]
  assign io_sigs_fma = _T_81 | decoder_4; // @[FPU.scala 133:40]
  assign io_sigs_div = _T_82 == 32'h18000010; // @[FPU.scala 133:40]
  assign io_sigs_sqrt = _T_73 == 32'h50000010; // @[FPU.scala 133:40]
  assign io_sigs_wflags = _T_94 | _T_91; // @[FPU.scala 133:40]
  assign FPUDecoder_covSum = 30'h0;
  assign io_covSum = FPUDecoder_covSum;
  assign metaAssert = 1'h0;
endmodule
module FPUFMAPipe(
  input         clock,
  input         reset,
  input         io_in_valid,
  input         io_in_bits_ren3,
  input         io_in_bits_swap23,
  input  [2:0]  io_in_bits_rm,
  input  [1:0]  io_in_bits_fmaCmd,
  input  [64:0] io_in_bits_in1,
  input  [64:0] io_in_bits_in2,
  input  [64:0] io_in_bits_in3,
  output [64:0] io_out_bits_data,
  output [4:0]  io_out_bits_exc,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         fma_halt
);
  wire  fma_clock; // @[FPU.scala 644:19]
  wire  fma_reset; // @[FPU.scala 644:19]
  wire  fma_io_validin; // @[FPU.scala 644:19]
  wire [1:0] fma_io_op; // @[FPU.scala 644:19]
  wire [32:0] fma_io_a; // @[FPU.scala 644:19]
  wire [32:0] fma_io_b; // @[FPU.scala 644:19]
  wire [32:0] fma_io_c; // @[FPU.scala 644:19]
  wire [2:0] fma_io_roundingMode; // @[FPU.scala 644:19]
  wire [32:0] fma_io_out; // @[FPU.scala 644:19]
  wire [4:0] fma_io_exceptionFlags; // @[FPU.scala 644:19]
  wire [29:0] fma_io_covSum; // @[FPU.scala 644:19]
  wire  fma_metaAssert; // @[FPU.scala 644:19]
  wire  fma_metaReset; // @[FPU.scala 644:19]
  reg  valid; // @[FPU.scala 632:18]
  reg [31:0] _RAND_0;
  reg [2:0] in_rm; // @[FPU.scala 633:15]
  reg [31:0] _RAND_1;
  reg [1:0] in_fmaCmd; // @[FPU.scala 633:15]
  reg [31:0] _RAND_2;
  reg [64:0] in_in1; // @[FPU.scala 633:15]
  reg [95:0] _RAND_3;
  reg [64:0] in_in2; // @[FPU.scala 633:15]
  reg [95:0] _RAND_4;
  reg [64:0] in_in3; // @[FPU.scala 633:15]
  reg [95:0] _RAND_5;
  wire [64:0] _T_13; // @[FPU.scala 636:32]
  wire [64:0] _T_15; // @[FPU.scala 636:50]
  wire  _T_16; // @[FPU.scala 641:21]
  wire [29:0] FPUFMAPipe_covSum;
  wire [29:0] fma_sum;
  wire  fma_metaAssert_wire;
  reg  FPUFMAPipe_metaAssert;
  reg [31:0] _RAND_6;
  MulAddRecFNPipe fma ( // @[FPU.scala 644:19]
    .clock(fma_clock),
    .reset(fma_reset),
    .io_validin(fma_io_validin),
    .io_op(fma_io_op),
    .io_a(fma_io_a),
    .io_b(fma_io_b),
    .io_c(fma_io_c),
    .io_roundingMode(fma_io_roundingMode),
    .io_out(fma_io_out),
    .io_exceptionFlags(fma_io_exceptionFlags),
    .io_covSum(fma_io_covSum),
    .metaAssert(fma_metaAssert),
    .metaReset(fma_metaReset)
  );
  assign _T_13 = io_in_bits_in1 ^ io_in_bits_in2; // @[FPU.scala 636:32]
  assign _T_15 = _T_13 & 65'h100000000; // @[FPU.scala 636:50]
  assign _T_16 = io_in_bits_ren3 | io_in_bits_swap23; // @[FPU.scala 641:21]
  assign io_out_bits_data = {{32'd0}, fma_io_out}; // @[FPU.scala 657:10]
  assign io_out_bits_exc = fma_io_exceptionFlags; // @[FPU.scala 657:10]
  assign fma_clock = clock;
  assign fma_reset = reset;
  assign fma_io_validin = valid; // @[FPU.scala 645:18]
  assign fma_io_op = in_fmaCmd; // @[FPU.scala 646:13]
  assign fma_io_a = in_in1[32:0]; // @[FPU.scala 649:12]
  assign fma_io_b = in_in2[32:0]; // @[FPU.scala 650:12]
  assign fma_io_c = in_in3[32:0]; // @[FPU.scala 651:12]
  assign fma_io_roundingMode = in_rm; // @[FPU.scala 647:23]
  assign FPUFMAPipe_covSum = 30'h0;
  assign fma_sum = FPUFMAPipe_covSum + fma_io_covSum;
  assign io_covSum = fma_sum;
  assign fma_metaAssert_wire = fma_metaAssert;
  assign metaAssert = FPUFMAPipe_metaAssert;
  assign fma_metaReset = metaReset | fma_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_rm = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_fmaCmd = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {3{`RANDOM}};
  in_in1 = _RAND_3[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {3{`RANDOM}};
  in_in2 = _RAND_4[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {3{`RANDOM}};
  in_in3 = _RAND_5[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  FPUFMAPipe_metaAssert = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      valid <= 1'h0;
    end else begin
      valid <= io_in_valid;
    end
    if (metaReset) begin
      in_rm <= 3'h0;
    end else if (io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if (metaReset) begin
      in_fmaCmd <= 2'h0;
    end else if (io_in_valid) begin
      in_fmaCmd <= io_in_bits_fmaCmd;
    end
    if (metaReset) begin
      in_in1 <= 65'h0;
    end else if (io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if (metaReset) begin
      in_in2 <= 65'h0;
    end else if (io_in_valid) begin
      if (io_in_bits_swap23) begin
        in_in2 <= 65'h80000000;
      end else begin
        in_in2 <= io_in_bits_in2;
      end
    end
    if (metaReset) begin
      in_in3 <= 65'h0;
    end else if (io_in_valid) begin
      if (~_T_16) begin
        in_in3 <= _T_15;
      end else begin
        in_in3 <= io_in_bits_in3;
      end
    end
    if (metaReset) begin
      FPUFMAPipe_metaAssert <= 1'h0;
    end else begin
      FPUFMAPipe_metaAssert <= FPUFMAPipe_metaAssert | fma_metaAssert_wire;
    end
  end
endmodule
module FPToInt(
  input         clock,
  input         io_in_valid,
  input         io_in_bits_ren2,
  input         io_in_bits_singleIn,
  input         io_in_bits_singleOut,
  input         io_in_bits_wflags,
  input  [2:0]  io_in_bits_rm,
  input  [1:0]  io_in_bits_typ,
  input  [64:0] io_in_bits_in1,
  input  [64:0] io_in_bits_in2,
  output [2:0]  io_out_bits_in_rm,
  output [64:0] io_out_bits_in_in1,
  output [64:0] io_out_bits_in_in2,
  output        io_out_bits_lt,
  output [63:0] io_out_bits_store,
  output [63:0] io_out_bits_toint,
  output [4:0]  io_out_bits_exc,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [64:0] dcmp_io_a; // @[FPU.scala 397:20]
  wire [64:0] dcmp_io_b; // @[FPU.scala 397:20]
  wire  dcmp_io_signaling; // @[FPU.scala 397:20]
  wire  dcmp_io_lt; // @[FPU.scala 397:20]
  wire  dcmp_io_eq; // @[FPU.scala 397:20]
  wire [4:0] dcmp_io_exceptionFlags; // @[FPU.scala 397:20]
  wire [29:0] dcmp_io_covSum; // @[FPU.scala 397:20]
  wire  dcmp_metaAssert; // @[FPU.scala 397:20]
  wire [64:0] RecFNToIN_io_in; // @[FPU.scala 425:24]
  wire [2:0] RecFNToIN_io_roundingMode; // @[FPU.scala 425:24]
  wire  RecFNToIN_io_signedOut; // @[FPU.scala 425:24]
  wire [63:0] RecFNToIN_io_out; // @[FPU.scala 425:24]
  wire [2:0] RecFNToIN_io_intExceptionFlags; // @[FPU.scala 425:24]
  wire [29:0] RecFNToIN_io_covSum; // @[FPU.scala 425:24]
  wire  RecFNToIN_metaAssert; // @[FPU.scala 425:24]
  wire [64:0] RecFNToIN_1_io_in; // @[FPU.scala 435:30]
  wire [2:0] RecFNToIN_1_io_roundingMode; // @[FPU.scala 435:30]
  wire  RecFNToIN_1_io_signedOut; // @[FPU.scala 435:30]
  wire [2:0] RecFNToIN_1_io_intExceptionFlags; // @[FPU.scala 435:30]
  wire [29:0] RecFNToIN_1_io_covSum; // @[FPU.scala 435:30]
  wire  RecFNToIN_1_metaAssert; // @[FPU.scala 435:30]
  reg  in_ren2; // @[Reg.scala 11:16]
  reg [31:0] _RAND_0;
  reg  in_singleOut; // @[Reg.scala 11:16]
  reg [31:0] _RAND_1;
  reg  in_wflags; // @[Reg.scala 11:16]
  reg [31:0] _RAND_2;
  reg [2:0] in_rm; // @[Reg.scala 11:16]
  reg [31:0] _RAND_3;
  reg [1:0] in_typ; // @[Reg.scala 11:16]
  reg [31:0] _RAND_4;
  reg [64:0] in_in1; // @[Reg.scala 11:16]
  reg [95:0] _RAND_5;
  reg [64:0] in_in2; // @[Reg.scala 11:16]
  reg [95:0] _RAND_6;
  wire  tag; // @[FPU.scala 402:13]
  wire  _T_16; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_18; // @[rawFloatFromRecFN.scala 52:54]
  wire  _T_22; // @[rawFloatFromRecFN.scala 55:33]
  wire  _T_25; // @[rawFloatFromRecFN.scala 56:33]
  wire [12:0] _T_27; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] _T_31; // @[Cat.scala 30:58]
  wire  _T_32; // @[fNFromRecFN.scala 50:39]
  wire [5:0] _T_36; // @[fNFromRecFN.scala 51:39]
  wire [52:0] _T_38; // @[fNFromRecFN.scala 52:42]
  wire [10:0] _T_43; // @[fNFromRecFN.scala 57:45]
  wire [10:0] _T_44; // @[fNFromRecFN.scala 55:16]
  wire  _T_45; // @[fNFromRecFN.scala 59:44]
  wire [10:0] _T_47; // @[Bitwise.scala 72:12]
  wire [10:0] _T_48; // @[fNFromRecFN.scala 59:15]
  wire [51:0] _T_50; // @[fNFromRecFN.scala 63:20]
  wire [51:0] _T_51; // @[fNFromRecFN.scala 61:16]
  wire [63:0] _T_53; // @[Cat.scala 30:58]
  wire [32:0] _T_58; // @[Cat.scala 30:58]
  wire  _T_61; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_63; // @[rawFloatFromRecFN.scala 52:54]
  wire  _T_67; // @[rawFloatFromRecFN.scala 55:33]
  wire  _T_70; // @[rawFloatFromRecFN.scala 56:33]
  wire [9:0] _T_72; // @[rawFloatFromRecFN.scala 59:27]
  wire [24:0] _T_76; // @[Cat.scala 30:58]
  wire  _T_77; // @[fNFromRecFN.scala 50:39]
  wire [4:0] _T_81; // @[fNFromRecFN.scala 51:39]
  wire [23:0] _T_83; // @[fNFromRecFN.scala 52:42]
  wire [7:0] _T_88; // @[fNFromRecFN.scala 57:45]
  wire [7:0] _T_89; // @[fNFromRecFN.scala 55:16]
  wire  _T_90; // @[fNFromRecFN.scala 59:44]
  wire [7:0] _T_92; // @[Bitwise.scala 72:12]
  wire [7:0] _T_93; // @[fNFromRecFN.scala 59:15]
  wire [22:0] _T_95; // @[fNFromRecFN.scala 63:20]
  wire [22:0] _T_96; // @[fNFromRecFN.scala 61:16]
  wire [31:0] _T_98; // @[Cat.scala 30:58]
  wire  _T_102; // @[FPU.scala 197:56]
  wire [31:0] _T_104; // @[FPU.scala 373:44]
  wire [63:0] store; // @[Cat.scala 30:58]
  wire [63:0] _T_108; // @[Cat.scala 30:58]
  wire  _T_272; // @[FPU.scala 442:54]
  wire  _T_264; // @[FPU.scala 440:59]
  wire  _T_265; // @[FPU.scala 441:46]
  wire [30:0] _T_268; // @[Bitwise.scala 72:12]
  wire [63:0] _T_274; // @[Cat.scala 30:58]
  wire [63:0] _GEN_24; // @[FPU.scala 443:26]
  wire [63:0] _GEN_25; // @[FPU.scala 434:30]
  wire [1:0] _T_241; // @[Cat.scala 30:58]
  wire [2:0] _GEN_33; // @[FPU.scala 417:22]
  wire [2:0] _T_242; // @[FPU.scala 417:22]
  wire  _T_243; // @[FPU.scala 417:53]
  wire [63:0] _T_245; // @[FPU.scala 417:77]
  wire [63:0] _GEN_34; // @[FPU.scala 417:57]
  wire [63:0] _T_246; // @[FPU.scala 417:57]
  wire [63:0] _GEN_28; // @[FPU.scala 421:21]
  wire  _T_213; // @[FPU.scala 213:24]
  wire  _T_211; // @[FPU.scala 212:24]
  wire  _T_191; // @[FPU.scala 204:28]
  wire  _T_206; // @[FPU.scala 210:27]
  wire  _T_215; // @[FPU.scala 215:31]
  wire  _T_198; // @[FPU.scala 208:27]
  wire  _T_193; // @[FPU.scala 206:55]
  wire  _T_200; // @[FPU.scala 208:39]
  wire  _T_201; // @[FPU.scala 208:71]
  wire  _T_202; // @[FPU.scala 208:61]
  wire  _T_217; // @[FPU.scala 215:50]
  wire  _T_194; // @[FPU.scala 207:28]
  wire  _T_196; // @[FPU.scala 207:62]
  wire  _T_197; // @[FPU.scala 207:40]
  wire  _T_219; // @[FPU.scala 216:21]
  wire  _T_203; // @[FPU.scala 209:23]
  wire  _T_221; // @[FPU.scala 216:38]
  wire  _T_222; // @[FPU.scala 216:55]
  wire  _T_223; // @[FPU.scala 217:21]
  wire  _T_224; // @[FPU.scala 217:39]
  wire  _T_225; // @[FPU.scala 217:54]
  wire [9:0] _T_234; // @[Cat.scala 30:58]
  wire  _T_133; // @[FPU.scala 229:36]
  wire  _T_134; // @[FPU.scala 229:25]
  wire [11:0] _T_128; // @[FPU.scala 228:31]
  wire [11:0] _T_131; // @[FPU.scala 228:48]
  wire [8:0] _T_136; // @[Cat.scala 30:58]
  wire [8:0] _T_138; // @[FPU.scala 229:10]
  wire [75:0] _T_124; // @[FPU.scala 225:28]
  wire [32:0] _T_140; // @[Cat.scala 30:58]
  wire  _T_161; // @[FPU.scala 211:22]
  wire  _T_166; // @[FPU.scala 213:24]
  wire  _T_164; // @[FPU.scala 212:24]
  wire  _T_144; // @[FPU.scala 204:28]
  wire  _T_159; // @[FPU.scala 210:27]
  wire  _T_168; // @[FPU.scala 215:31]
  wire  _T_151; // @[FPU.scala 208:27]
  wire  _T_146; // @[FPU.scala 206:55]
  wire  _T_153; // @[FPU.scala 208:39]
  wire  _T_154; // @[FPU.scala 208:71]
  wire  _T_155; // @[FPU.scala 208:61]
  wire  _T_170; // @[FPU.scala 215:50]
  wire  _T_147; // @[FPU.scala 207:28]
  wire  _T_149; // @[FPU.scala 207:62]
  wire  _T_150; // @[FPU.scala 207:40]
  wire  _T_172; // @[FPU.scala 216:21]
  wire  _T_156; // @[FPU.scala 209:23]
  wire  _T_174; // @[FPU.scala 216:38]
  wire  _T_175; // @[FPU.scala 216:55]
  wire  _T_176; // @[FPU.scala 217:21]
  wire  _T_177; // @[FPU.scala 217:39]
  wire  _T_178; // @[FPU.scala 217:54]
  wire [9:0] _T_187; // @[Cat.scala 30:58]
  wire [9:0] _T_236; // @[package.scala 31:71]
  wire [63:0] _GEN_35; // @[FPU.scala 412:27]
  wire [63:0] _T_239; // @[FPU.scala 412:27]
  wire [63:0] _GEN_22; // @[FPU.scala 410:19]
  wire [63:0] toint; // @[FPU.scala 416:20]
  wire [31:0] _T_115; // @[Bitwise.scala 72:12]
  wire [63:0] _T_116; // @[Cat.scala 30:58]
  wire  _GEN_27; // @[FPU.scala 421:21]
  wire  _GEN_23; // @[FPU.scala 410:19]
  wire  intType; // @[FPU.scala 416:20]
  wire  _T_252; // @[FPU.scala 430:62]
  wire [4:0] _T_255; // @[Cat.scala 30:58]
  wire  _T_277; // @[FPU.scala 444:64]
  wire [4:0] _T_279; // @[Cat.scala 30:58]
  wire [4:0] _GEN_26; // @[FPU.scala 434:30]
  wire [4:0] _GEN_29; // @[FPU.scala 421:21]
  wire  _T_281; // @[FPU.scala 451:53]
  wire  _T_283; // @[FPU.scala 451:79]
  wire  _T_284; // @[FPU.scala 451:59]
  reg [4:0] FPToInt_state; // @[Register tracking FPToInt state]
  reg [31:0] _RAND_7;
  reg  FPToInt_cov [0:31]; // @[Coverage map for FPToInt]
  reg [31:0] _RAND_8;
  wire  FPToInt_cov_read_data; // @[Coverage map for FPToInt]
  wire [4:0] FPToInt_cov_read_addr; // @[Coverage map for FPToInt]
  wire  FPToInt_cov_write_data; // @[Coverage map for FPToInt]
  wire [4:0] FPToInt_cov_write_addr; // @[Coverage map for FPToInt]
  wire  FPToInt_cov_write_mask; // @[Coverage map for FPToInt]
  wire  FPToInt_cov_write_en; // @[Coverage map for FPToInt]
  reg [29:0] FPToInt_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_9;
  wire [1:0] in_typ_shl;
  wire [4:0] in_typ_pad;
  wire [2:0] in_singleOut_shl;
  wire [4:0] in_singleOut_pad;
  wire [3:0] in_ren2_shl;
  wire [4:0] in_ren2_pad;
  wire [4:0] in_wflags_shl;
  wire [4:0] in_wflags_pad;
  wire [4:0] FPToInt_xor1;
  wire [4:0] FPToInt_xor2;
  wire [4:0] FPToInt_xor0;
  wire [29:0] dcmp_sum;
  wire [29:0] RecFNToIN_sum;
  wire [29:0] RecFNToIN_1_sum;
  wire  dcmp_metaAssert_wire;
  wire  RecFNToIN_metaAssert_wire;
  wire  RecFNToIN_1_metaAssert_wire;
  wire  FPToInt_or2;
  wire  FPToInt_or0;
  CompareRecFN dcmp ( // @[FPU.scala 397:20]
    .io_a(dcmp_io_a),
    .io_b(dcmp_io_b),
    .io_signaling(dcmp_io_signaling),
    .io_lt(dcmp_io_lt),
    .io_eq(dcmp_io_eq),
    .io_exceptionFlags(dcmp_io_exceptionFlags),
    .io_covSum(dcmp_io_covSum),
    .metaAssert(dcmp_metaAssert)
  );
  RecFNToIN RecFNToIN ( // @[FPU.scala 425:24]
    .io_in(RecFNToIN_io_in),
    .io_roundingMode(RecFNToIN_io_roundingMode),
    .io_signedOut(RecFNToIN_io_signedOut),
    .io_out(RecFNToIN_io_out),
    .io_intExceptionFlags(RecFNToIN_io_intExceptionFlags),
    .io_covSum(RecFNToIN_io_covSum),
    .metaAssert(RecFNToIN_metaAssert)
  );
  RecFNToIN_1 RecFNToIN_1 ( // @[FPU.scala 435:30]
    .io_in(RecFNToIN_1_io_in),
    .io_roundingMode(RecFNToIN_1_io_roundingMode),
    .io_signedOut(RecFNToIN_1_io_signedOut),
    .io_intExceptionFlags(RecFNToIN_1_io_intExceptionFlags),
    .io_covSum(RecFNToIN_1_io_covSum),
    .metaAssert(RecFNToIN_1_metaAssert)
  );
  assign tag = ~in_singleOut; // @[FPU.scala 402:13]
  assign _T_16 = in_in1[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_18 = in_in1[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign _T_22 = _T_18 & in_in1[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign _T_25 = _T_18 & ~in_in1[61]; // @[rawFloatFromRecFN.scala 56:33]
  assign _T_27 = {1'b0,$signed(in_in1[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign _T_31 = {1'h0,~_T_16,in_in1[51:0]}; // @[Cat.scala 30:58]
  assign _T_32 = $signed(_T_27) < 13'sh402; // @[fNFromRecFN.scala 50:39]
  assign _T_36 = 6'h1 - _T_27[5:0]; // @[fNFromRecFN.scala 51:39]
  assign _T_38 = _T_31[53:1] >> _T_36; // @[fNFromRecFN.scala 52:42]
  assign _T_43 = _T_27[10:0] - 11'h401; // @[fNFromRecFN.scala 57:45]
  assign _T_44 = _T_32 ? 11'h0 : _T_43; // @[fNFromRecFN.scala 55:16]
  assign _T_45 = _T_22 | _T_25; // @[fNFromRecFN.scala 59:44]
  assign _T_47 = _T_45 ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  assign _T_48 = _T_44 | _T_47; // @[fNFromRecFN.scala 59:15]
  assign _T_50 = _T_25 ? 52'h0 : _T_31[51:0]; // @[fNFromRecFN.scala 63:20]
  assign _T_51 = _T_32 ? _T_38[51:0] : _T_50; // @[fNFromRecFN.scala 61:16]
  assign _T_53 = {in_in1[64],_T_48,_T_51}; // @[Cat.scala 30:58]
  assign _T_58 = {in_in1[31],in_in1[52],in_in1[30:0]}; // @[Cat.scala 30:58]
  assign _T_61 = _T_58[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_63 = _T_58[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign _T_67 = _T_63 & _T_58[29]; // @[rawFloatFromRecFN.scala 55:33]
  assign _T_70 = _T_63 & ~_T_58[29]; // @[rawFloatFromRecFN.scala 56:33]
  assign _T_72 = {1'b0,$signed(_T_58[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  assign _T_76 = {1'h0,~_T_61,_T_58[22:0]}; // @[Cat.scala 30:58]
  assign _T_77 = $signed(_T_72) < 10'sh82; // @[fNFromRecFN.scala 50:39]
  assign _T_81 = 5'h1 - _T_72[4:0]; // @[fNFromRecFN.scala 51:39]
  assign _T_83 = _T_76[24:1] >> _T_81; // @[fNFromRecFN.scala 52:42]
  assign _T_88 = _T_72[7:0] - 8'h81; // @[fNFromRecFN.scala 57:45]
  assign _T_89 = _T_77 ? 8'h0 : _T_88; // @[fNFromRecFN.scala 55:16]
  assign _T_90 = _T_67 | _T_70; // @[fNFromRecFN.scala 59:44]
  assign _T_92 = _T_90 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_93 = _T_89 | _T_92; // @[fNFromRecFN.scala 59:15]
  assign _T_95 = _T_70 ? 23'h0 : _T_76[22:0]; // @[fNFromRecFN.scala 63:20]
  assign _T_96 = _T_77 ? _T_83[22:0] : _T_95; // @[fNFromRecFN.scala 61:16]
  assign _T_98 = {_T_58[32],_T_93,_T_96}; // @[Cat.scala 30:58]
  assign _T_102 = ~in_in1[63:61] == 3'h0; // @[FPU.scala 197:56]
  assign _T_104 = _T_102 ? _T_98 : _T_53[31:0]; // @[FPU.scala 373:44]
  assign store = {_T_53[63:32],_T_104}; // @[Cat.scala 30:58]
  assign _T_108 = {store[31:0],store[31:0]}; // @[Cat.scala 30:58]
  assign _T_272 = RecFNToIN_io_intExceptionFlags[2] | RecFNToIN_1_io_intExceptionFlags[1]; // @[FPU.scala 442:54]
  assign _T_264 = in_in1[64] & ~_T_102; // @[FPU.scala 440:59]
  assign _T_265 = RecFNToIN_io_signedOut == _T_264; // @[FPU.scala 441:46]
  assign _T_268 = _T_264 ? 31'h0 : 31'h7fffffff; // @[Bitwise.scala 72:12]
  assign _T_274 = {RecFNToIN_io_out[63:32],_T_265,_T_268}; // @[Cat.scala 30:58]
  assign _GEN_24 = _T_272 ? _T_274 : RecFNToIN_io_out; // @[FPU.scala 443:26]
  assign _GEN_25 = in_typ[1] ? RecFNToIN_io_out : _GEN_24; // @[FPU.scala 434:30]
  assign _T_241 = {dcmp_io_lt,dcmp_io_eq}; // @[Cat.scala 30:58]
  assign _GEN_33 = {{1'd0}, _T_241}; // @[FPU.scala 417:22]
  assign _T_242 = ~in_rm & _GEN_33; // @[FPU.scala 417:22]
  assign _T_243 = _T_242 != 3'h0; // @[FPU.scala 417:53]
  assign _T_245 = {store[63:32], 32'h0}; // @[FPU.scala 417:77]
  assign _GEN_34 = {{63'd0}, _T_243}; // @[FPU.scala 417:57]
  assign _T_246 = _GEN_34 | _T_245; // @[FPU.scala 417:57]
  assign _GEN_28 = in_ren2 ? _T_246 : _GEN_25; // @[FPU.scala 421:21]
  assign _T_213 = _T_102 & in_in1[51]; // @[FPU.scala 213:24]
  assign _T_211 = _T_102 & ~in_in1[51]; // @[FPU.scala 212:24]
  assign _T_191 = in_in1[63:62] == 2'h3; // @[FPU.scala 204:28]
  assign _T_206 = _T_191 & ~in_in1[61]; // @[FPU.scala 210:27]
  assign _T_215 = _T_206 & ~in_in1[64]; // @[FPU.scala 215:31]
  assign _T_198 = in_in1[63:62] == 2'h1; // @[FPU.scala 208:27]
  assign _T_193 = in_in1[61:52] < 10'h2; // @[FPU.scala 206:55]
  assign _T_200 = _T_198 & ~_T_193; // @[FPU.scala 208:39]
  assign _T_201 = in_in1[63:62] == 2'h2; // @[FPU.scala 208:71]
  assign _T_202 = _T_200 | _T_201; // @[FPU.scala 208:61]
  assign _T_217 = _T_202 & ~in_in1[64]; // @[FPU.scala 215:50]
  assign _T_194 = in_in1[63:61] == 3'h1; // @[FPU.scala 207:28]
  assign _T_196 = _T_198 & _T_193; // @[FPU.scala 207:62]
  assign _T_197 = _T_194 | _T_196; // @[FPU.scala 207:40]
  assign _T_219 = _T_197 & ~in_in1[64]; // @[FPU.scala 216:21]
  assign _T_203 = in_in1[63:61] == 3'h0; // @[FPU.scala 209:23]
  assign _T_221 = _T_203 & ~in_in1[64]; // @[FPU.scala 216:38]
  assign _T_222 = _T_203 & in_in1[64]; // @[FPU.scala 216:55]
  assign _T_223 = _T_197 & in_in1[64]; // @[FPU.scala 217:21]
  assign _T_224 = _T_202 & in_in1[64]; // @[FPU.scala 217:39]
  assign _T_225 = _T_206 & in_in1[64]; // @[FPU.scala 217:54]
  assign _T_234 = {_T_213,_T_211,_T_215,_T_217,_T_219,_T_221,_T_222,_T_223,_T_224,_T_225}; // @[Cat.scala 30:58]
  assign _T_133 = in_in1[63:61] >= 3'h6; // @[FPU.scala 229:36]
  assign _T_134 = _T_16 | _T_133; // @[FPU.scala 229:25]
  assign _T_128 = in_in1[63:52] + 12'h100; // @[FPU.scala 228:31]
  assign _T_131 = _T_128 - 12'h800; // @[FPU.scala 228:48]
  assign _T_136 = {in_in1[63:61],_T_131[5:0]}; // @[Cat.scala 30:58]
  assign _T_138 = _T_134 ? _T_136 : _T_131[8:0]; // @[FPU.scala 229:10]
  assign _T_124 = {in_in1[51:0], 24'h0}; // @[FPU.scala 225:28]
  assign _T_140 = {in_in1[64],_T_138,_T_124[75:53]}; // @[Cat.scala 30:58]
  assign _T_161 = ~_T_140[31:29] == 3'h0; // @[FPU.scala 211:22]
  assign _T_166 = _T_161 & _T_140[22]; // @[FPU.scala 213:24]
  assign _T_164 = _T_161 & ~_T_140[22]; // @[FPU.scala 212:24]
  assign _T_144 = _T_140[31:30] == 2'h3; // @[FPU.scala 204:28]
  assign _T_159 = _T_144 & ~_T_140[29]; // @[FPU.scala 210:27]
  assign _T_168 = _T_159 & ~_T_140[32]; // @[FPU.scala 215:31]
  assign _T_151 = _T_140[31:30] == 2'h1; // @[FPU.scala 208:27]
  assign _T_146 = _T_140[29:23] < 7'h2; // @[FPU.scala 206:55]
  assign _T_153 = _T_151 & ~_T_146; // @[FPU.scala 208:39]
  assign _T_154 = _T_140[31:30] == 2'h2; // @[FPU.scala 208:71]
  assign _T_155 = _T_153 | _T_154; // @[FPU.scala 208:61]
  assign _T_170 = _T_155 & ~_T_140[32]; // @[FPU.scala 215:50]
  assign _T_147 = _T_140[31:29] == 3'h1; // @[FPU.scala 207:28]
  assign _T_149 = _T_151 & _T_146; // @[FPU.scala 207:62]
  assign _T_150 = _T_147 | _T_149; // @[FPU.scala 207:40]
  assign _T_172 = _T_150 & ~_T_140[32]; // @[FPU.scala 216:21]
  assign _T_156 = _T_140[31:29] == 3'h0; // @[FPU.scala 209:23]
  assign _T_174 = _T_156 & ~_T_140[32]; // @[FPU.scala 216:38]
  assign _T_175 = _T_156 & _T_140[32]; // @[FPU.scala 216:55]
  assign _T_176 = _T_150 & _T_140[32]; // @[FPU.scala 217:21]
  assign _T_177 = _T_155 & _T_140[32]; // @[FPU.scala 217:39]
  assign _T_178 = _T_159 & _T_140[32]; // @[FPU.scala 217:54]
  assign _T_187 = {_T_166,_T_164,_T_168,_T_170,_T_172,_T_174,_T_175,_T_176,_T_177,_T_178}; // @[Cat.scala 30:58]
  assign _T_236 = tag ? _T_234 : _T_187; // @[package.scala 31:71]
  assign _GEN_35 = {{54'd0}, _T_236}; // @[FPU.scala 412:27]
  assign _T_239 = _GEN_35 | _T_245; // @[FPU.scala 412:27]
  assign _GEN_22 = in_rm[0] ? _T_239 : store; // @[FPU.scala 410:19]
  assign toint = in_wflags ? _GEN_28 : _GEN_22; // @[FPU.scala 416:20]
  assign _T_115 = toint[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  assign _T_116 = {_T_115,toint[31:0]}; // @[Cat.scala 30:58]
  assign _GEN_27 = ~in_ren2 & in_typ[1]; // @[FPU.scala 421:21]
  assign _GEN_23 = in_rm[0] ? 1'h0 : tag; // @[FPU.scala 410:19]
  assign intType = in_wflags ? _GEN_27 : _GEN_23; // @[FPU.scala 416:20]
  assign _T_252 = RecFNToIN_io_intExceptionFlags[2:1] != 2'h0; // @[FPU.scala 430:62]
  assign _T_255 = {_T_252,3'h0,RecFNToIN_io_intExceptionFlags[0]}; // @[Cat.scala 30:58]
  assign _T_277 = ~_T_272 & RecFNToIN_io_intExceptionFlags[0]; // @[FPU.scala 444:64]
  assign _T_279 = {_T_272,3'h0,_T_277}; // @[Cat.scala 30:58]
  assign _GEN_26 = in_typ[1] ? _T_255 : _T_279; // @[FPU.scala 434:30]
  assign _GEN_29 = in_ren2 ? dcmp_io_exceptionFlags : _GEN_26; // @[FPU.scala 421:21]
  assign _T_281 = $signed(dcmp_io_a) < 65'sh0; // @[FPU.scala 451:53]
  assign _T_283 = $signed(dcmp_io_b) >= 65'sh0; // @[FPU.scala 451:79]
  assign _T_284 = _T_281 & _T_283; // @[FPU.scala 451:59]
  assign io_out_bits_in_rm = in_rm; // @[FPU.scala 452:18]
  assign io_out_bits_in_in1 = in_in1; // @[FPU.scala 452:18]
  assign io_out_bits_in_in2 = in_in2; // @[FPU.scala 452:18]
  assign io_out_bits_lt = dcmp_io_lt | _T_284; // @[FPU.scala 451:18]
  assign io_out_bits_store = tag ? store : _T_108; // @[FPU.scala 406:21]
  assign io_out_bits_toint = intType ? toint : _T_116; // @[FPU.scala 407:21]
  assign io_out_bits_exc = in_wflags ? _GEN_29 : 5'h0; // @[FPU.scala 408:19 FPU.scala 418:21 FPU.scala 430:23 FPU.scala 444:27]
  assign dcmp_io_a = in_in1; // @[FPU.scala 398:13]
  assign dcmp_io_b = in_in2; // @[FPU.scala 399:13]
  assign dcmp_io_signaling = ~in_rm[1]; // @[FPU.scala 400:21]
  assign RecFNToIN_io_in = in_in1; // @[FPU.scala 426:18]
  assign RecFNToIN_io_roundingMode = in_rm; // @[FPU.scala 427:28]
  assign RecFNToIN_io_signedOut = ~in_typ[0]; // @[FPU.scala 428:25]
  assign RecFNToIN_1_io_in = in_in1; // @[FPU.scala 436:24]
  assign RecFNToIN_1_io_roundingMode = in_rm; // @[FPU.scala 437:34]
  assign RecFNToIN_1_io_signedOut = ~in_typ[0]; // @[FPU.scala 438:31]
  assign FPToInt_cov_read_addr = FPToInt_state;
  assign FPToInt_cov_read_data = FPToInt_cov[FPToInt_cov_read_addr]; // @[Coverage map for FPToInt]
  assign FPToInt_cov_write_data = 1'h1;
  assign FPToInt_cov_write_addr = FPToInt_state;
  assign FPToInt_cov_write_mask = 1'h1;
  assign FPToInt_cov_write_en = 1'h1;
  assign in_typ_shl = in_typ;
  assign in_typ_pad = {3'h0,in_typ_shl};
  assign in_singleOut_shl = {in_singleOut, 2'h0};
  assign in_singleOut_pad = {2'h0,in_singleOut_shl};
  assign in_ren2_shl = {in_ren2, 3'h0};
  assign in_ren2_pad = {1'h0,in_ren2_shl};
  assign in_wflags_shl = {in_wflags, 4'h0};
  assign in_wflags_pad = in_wflags_shl;
  assign FPToInt_xor1 = in_typ_pad ^ in_singleOut_pad;
  assign FPToInt_xor2 = in_ren2_pad ^ in_wflags_pad;
  assign FPToInt_xor0 = FPToInt_xor1 ^ FPToInt_xor2;
  assign dcmp_sum = FPToInt_covSum + dcmp_io_covSum;
  assign RecFNToIN_sum = dcmp_sum + RecFNToIN_io_covSum;
  assign RecFNToIN_1_sum = RecFNToIN_sum + RecFNToIN_1_io_covSum;
  assign io_covSum = RecFNToIN_1_sum;
  assign dcmp_metaAssert_wire = dcmp_metaAssert;
  assign RecFNToIN_metaAssert_wire = RecFNToIN_metaAssert;
  assign RecFNToIN_1_metaAssert_wire = RecFNToIN_1_metaAssert;
  assign FPToInt_or2 = RecFNToIN_metaAssert_wire | RecFNToIN_1_metaAssert_wire;
  assign FPToInt_or0 = dcmp_metaAssert_wire | FPToInt_or2;
  assign metaAssert = FPToInt_or0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_ren2 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_singleOut = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_wflags = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_rm = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  in_typ = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {3{`RANDOM}};
  in_in1 = _RAND_5[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {3{`RANDOM}};
  in_in2 = _RAND_6[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  FPToInt_state = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    FPToInt_cov[initvar] = _RAND_8[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  FPToInt_covSum = _RAND_9[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      in_ren2 <= 1'h0;
    end else if (io_in_valid) begin
      in_ren2 <= io_in_bits_ren2;
    end
    if (metaReset) begin
      in_singleOut <= 1'h0;
    end else if (io_in_valid) begin
      in_singleOut <= io_in_bits_singleOut;
    end
    if (metaReset) begin
      in_wflags <= 1'h0;
    end else if (io_in_valid) begin
      in_wflags <= io_in_bits_wflags;
    end
    if (metaReset) begin
      in_rm <= 3'h0;
    end else if (io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if (metaReset) begin
      in_typ <= 2'h0;
    end else if (io_in_valid) begin
      in_typ <= io_in_bits_typ;
    end
    if (metaReset) begin
      in_in1 <= 65'h0;
    end else if (io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if (metaReset) begin
      in_in2 <= 65'h0;
    end else if (io_in_valid) begin
      in_in2 <= io_in_bits_in2;
    end
    FPToInt_state <= FPToInt_xor0;
    if (!(FPToInt_cov_read_data)) begin
      FPToInt_covSum <= FPToInt_covSum + 1'h1;
    end
  end
  always @(posedge clock) begin
    if(FPToInt_cov_write_en & FPToInt_cov_write_mask) begin
      FPToInt_cov[FPToInt_cov_write_addr] <= FPToInt_cov_write_data; // @[Coverage map for FPToInt]
    end
  end
endmodule
module IntToFP(
  input         clock,
  input         reset,
  input         io_in_valid,
  input         io_in_bits_singleIn,
  input         io_in_bits_wflags,
  input  [2:0]  io_in_bits_rm,
  input  [1:0]  io_in_bits_typ,
  input  [63:0] io_in_bits_in1,
  output [64:0] io_out_bits_data,
  output [4:0]  io_out_bits_exc,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire  INToRecFN_io_signedIn; // @[FPU.scala 483:23]
  wire [63:0] INToRecFN_io_in; // @[FPU.scala 483:23]
  wire [2:0] INToRecFN_io_roundingMode; // @[FPU.scala 483:23]
  wire [32:0] INToRecFN_io_out; // @[FPU.scala 483:23]
  wire [4:0] INToRecFN_io_exceptionFlags; // @[FPU.scala 483:23]
  wire [29:0] INToRecFN_io_covSum; // @[FPU.scala 483:23]
  wire  INToRecFN_metaAssert; // @[FPU.scala 483:23]
  wire  INToRecFN_1_io_signedIn; // @[FPU.scala 483:23]
  wire [63:0] INToRecFN_1_io_in; // @[FPU.scala 483:23]
  wire [2:0] INToRecFN_1_io_roundingMode; // @[FPU.scala 483:23]
  wire [64:0] INToRecFN_1_io_out; // @[FPU.scala 483:23]
  wire [4:0] INToRecFN_1_io_exceptionFlags; // @[FPU.scala 483:23]
  wire [29:0] INToRecFN_1_io_covSum; // @[FPU.scala 483:23]
  wire  INToRecFN_1_metaAssert; // @[FPU.scala 483:23]
  reg  in_valid; // @[Valid.scala 48:22]
  reg [31:0] _RAND_0;
  reg  in_bits_singleIn; // @[Reg.scala 11:16]
  reg [31:0] _RAND_1;
  reg  in_bits_wflags; // @[Reg.scala 11:16]
  reg [31:0] _RAND_2;
  reg [2:0] in_bits_rm; // @[Reg.scala 11:16]
  reg [31:0] _RAND_3;
  reg [1:0] in_bits_typ; // @[Reg.scala 11:16]
  reg [31:0] _RAND_4;
  reg [63:0] in_bits_in1; // @[Reg.scala 11:16]
  reg [63:0] _RAND_5;
  wire  tag; // @[FPU.scala 462:13]
  wire [63:0] _T_21; // @[package.scala 31:71]
  wire [63:0] _T_22; // @[FPU.scala 358:23]
  wire  _T_26; // @[rawFloatFromFN.scala 50:34]
  wire  _T_27; // @[rawFloatFromFN.scala 51:38]
  wire [31:0] _T_32; // @[Bitwise.scala 103:31]
  wire [31:0] _T_34; // @[Bitwise.scala 103:65]
  wire [31:0] _T_36; // @[Bitwise.scala 103:75]
  wire [31:0] _T_37; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_24; // @[Bitwise.scala 103:31]
  wire [31:0] _T_42; // @[Bitwise.scala 103:31]
  wire [31:0] _T_44; // @[Bitwise.scala 103:65]
  wire [31:0] _T_46; // @[Bitwise.scala 103:75]
  wire [31:0] _T_47; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_25; // @[Bitwise.scala 103:31]
  wire [31:0] _T_52; // @[Bitwise.scala 103:31]
  wire [31:0] _T_54; // @[Bitwise.scala 103:65]
  wire [31:0] _T_56; // @[Bitwise.scala 103:75]
  wire [31:0] _T_57; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_26; // @[Bitwise.scala 103:31]
  wire [31:0] _T_62; // @[Bitwise.scala 103:31]
  wire [31:0] _T_64; // @[Bitwise.scala 103:65]
  wire [31:0] _T_66; // @[Bitwise.scala 103:75]
  wire [31:0] _T_67; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_27; // @[Bitwise.scala 103:31]
  wire [31:0] _T_72; // @[Bitwise.scala 103:31]
  wire [31:0] _T_74; // @[Bitwise.scala 103:65]
  wire [31:0] _T_76; // @[Bitwise.scala 103:75]
  wire [31:0] _T_77; // @[Bitwise.scala 103:39]
  wire [15:0] _T_83; // @[Bitwise.scala 103:31]
  wire [15:0] _T_85; // @[Bitwise.scala 103:65]
  wire [15:0] _T_87; // @[Bitwise.scala 103:75]
  wire [15:0] _T_88; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_28; // @[Bitwise.scala 103:31]
  wire [15:0] _T_93; // @[Bitwise.scala 103:31]
  wire [15:0] _T_95; // @[Bitwise.scala 103:65]
  wire [15:0] _T_97; // @[Bitwise.scala 103:75]
  wire [15:0] _T_98; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_29; // @[Bitwise.scala 103:31]
  wire [15:0] _T_103; // @[Bitwise.scala 103:31]
  wire [15:0] _T_105; // @[Bitwise.scala 103:65]
  wire [15:0] _T_107; // @[Bitwise.scala 103:75]
  wire [15:0] _T_108; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_30; // @[Bitwise.scala 103:31]
  wire [15:0] _T_113; // @[Bitwise.scala 103:31]
  wire [15:0] _T_115; // @[Bitwise.scala 103:65]
  wire [15:0] _T_117; // @[Bitwise.scala 103:75]
  wire [15:0] _T_118; // @[Bitwise.scala 103:39]
  wire [51:0] _T_130; // @[Cat.scala 30:58]
  wire [5:0] _T_183; // @[Mux.scala 31:69]
  wire [5:0] _T_184; // @[Mux.scala 31:69]
  wire [5:0] _T_185; // @[Mux.scala 31:69]
  wire [5:0] _T_186; // @[Mux.scala 31:69]
  wire [5:0] _T_187; // @[Mux.scala 31:69]
  wire [5:0] _T_188; // @[Mux.scala 31:69]
  wire [5:0] _T_189; // @[Mux.scala 31:69]
  wire [5:0] _T_190; // @[Mux.scala 31:69]
  wire [5:0] _T_191; // @[Mux.scala 31:69]
  wire [5:0] _T_192; // @[Mux.scala 31:69]
  wire [5:0] _T_193; // @[Mux.scala 31:69]
  wire [5:0] _T_194; // @[Mux.scala 31:69]
  wire [5:0] _T_195; // @[Mux.scala 31:69]
  wire [5:0] _T_196; // @[Mux.scala 31:69]
  wire [5:0] _T_197; // @[Mux.scala 31:69]
  wire [5:0] _T_198; // @[Mux.scala 31:69]
  wire [5:0] _T_199; // @[Mux.scala 31:69]
  wire [5:0] _T_200; // @[Mux.scala 31:69]
  wire [5:0] _T_201; // @[Mux.scala 31:69]
  wire [5:0] _T_202; // @[Mux.scala 31:69]
  wire [5:0] _T_203; // @[Mux.scala 31:69]
  wire [5:0] _T_204; // @[Mux.scala 31:69]
  wire [5:0] _T_205; // @[Mux.scala 31:69]
  wire [5:0] _T_206; // @[Mux.scala 31:69]
  wire [5:0] _T_207; // @[Mux.scala 31:69]
  wire [5:0] _T_208; // @[Mux.scala 31:69]
  wire [5:0] _T_209; // @[Mux.scala 31:69]
  wire [5:0] _T_210; // @[Mux.scala 31:69]
  wire [5:0] _T_211; // @[Mux.scala 31:69]
  wire [5:0] _T_212; // @[Mux.scala 31:69]
  wire [5:0] _T_213; // @[Mux.scala 31:69]
  wire [5:0] _T_214; // @[Mux.scala 31:69]
  wire [5:0] _T_215; // @[Mux.scala 31:69]
  wire [5:0] _T_216; // @[Mux.scala 31:69]
  wire [5:0] _T_217; // @[Mux.scala 31:69]
  wire [5:0] _T_218; // @[Mux.scala 31:69]
  wire [5:0] _T_219; // @[Mux.scala 31:69]
  wire [5:0] _T_220; // @[Mux.scala 31:69]
  wire [5:0] _T_221; // @[Mux.scala 31:69]
  wire [5:0] _T_222; // @[Mux.scala 31:69]
  wire [5:0] _T_223; // @[Mux.scala 31:69]
  wire [5:0] _T_224; // @[Mux.scala 31:69]
  wire [5:0] _T_225; // @[Mux.scala 31:69]
  wire [5:0] _T_226; // @[Mux.scala 31:69]
  wire [5:0] _T_227; // @[Mux.scala 31:69]
  wire [5:0] _T_228; // @[Mux.scala 31:69]
  wire [5:0] _T_229; // @[Mux.scala 31:69]
  wire [5:0] _T_230; // @[Mux.scala 31:69]
  wire [5:0] _T_231; // @[Mux.scala 31:69]
  wire [5:0] _T_232; // @[Mux.scala 31:69]
  wire [5:0] _T_233; // @[Mux.scala 31:69]
  wire [114:0] _GEN_31; // @[rawFloatFromFN.scala 54:36]
  wire [114:0] _T_234; // @[rawFloatFromFN.scala 54:36]
  wire [51:0] _T_236; // @[rawFloatFromFN.scala 54:64]
  wire [11:0] _GEN_32; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_237; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_238; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_239; // @[rawFloatFromFN.scala 60:27]
  wire [10:0] _GEN_33; // @[rawFloatFromFN.scala 60:22]
  wire [10:0] _T_240; // @[rawFloatFromFN.scala 60:22]
  wire [11:0] _GEN_34; // @[rawFloatFromFN.scala 59:15]
  wire [11:0] _T_242; // @[rawFloatFromFN.scala 59:15]
  wire  _T_243; // @[rawFloatFromFN.scala 62:34]
  wire  _T_245; // @[rawFloatFromFN.scala 63:62]
  wire  _T_249; // @[rawFloatFromFN.scala 66:33]
  wire [12:0] _T_252; // @[rawFloatFromFN.scala 70:48]
  wire [51:0] _T_254; // @[rawFloatFromFN.scala 72:42]
  wire [53:0] _T_256; // @[Cat.scala 30:58]
  wire [2:0] _T_258; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_35; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_260; // @[recFNFromFN.scala 48:79]
  wire [64:0] _T_265; // @[Cat.scala 30:58]
  wire  _T_269; // @[rawFloatFromFN.scala 50:34]
  wire  _T_270; // @[rawFloatFromFN.scala 51:38]
  wire [15:0] _T_275; // @[Bitwise.scala 103:31]
  wire [15:0] _T_277; // @[Bitwise.scala 103:65]
  wire [15:0] _T_279; // @[Bitwise.scala 103:75]
  wire [15:0] _T_280; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_36; // @[Bitwise.scala 103:31]
  wire [15:0] _T_285; // @[Bitwise.scala 103:31]
  wire [15:0] _T_287; // @[Bitwise.scala 103:65]
  wire [15:0] _T_289; // @[Bitwise.scala 103:75]
  wire [15:0] _T_290; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_37; // @[Bitwise.scala 103:31]
  wire [15:0] _T_295; // @[Bitwise.scala 103:31]
  wire [15:0] _T_297; // @[Bitwise.scala 103:65]
  wire [15:0] _T_299; // @[Bitwise.scala 103:75]
  wire [15:0] _T_300; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_38; // @[Bitwise.scala 103:31]
  wire [15:0] _T_305; // @[Bitwise.scala 103:31]
  wire [15:0] _T_307; // @[Bitwise.scala 103:65]
  wire [15:0] _T_309; // @[Bitwise.scala 103:75]
  wire [15:0] _T_310; // @[Bitwise.scala 103:39]
  wire [22:0] _T_330; // @[Cat.scala 30:58]
  wire [4:0] _T_354; // @[Mux.scala 31:69]
  wire [4:0] _T_355; // @[Mux.scala 31:69]
  wire [4:0] _T_356; // @[Mux.scala 31:69]
  wire [4:0] _T_357; // @[Mux.scala 31:69]
  wire [4:0] _T_358; // @[Mux.scala 31:69]
  wire [4:0] _T_359; // @[Mux.scala 31:69]
  wire [4:0] _T_360; // @[Mux.scala 31:69]
  wire [4:0] _T_361; // @[Mux.scala 31:69]
  wire [4:0] _T_362; // @[Mux.scala 31:69]
  wire [4:0] _T_363; // @[Mux.scala 31:69]
  wire [4:0] _T_364; // @[Mux.scala 31:69]
  wire [4:0] _T_365; // @[Mux.scala 31:69]
  wire [4:0] _T_366; // @[Mux.scala 31:69]
  wire [4:0] _T_367; // @[Mux.scala 31:69]
  wire [4:0] _T_368; // @[Mux.scala 31:69]
  wire [4:0] _T_369; // @[Mux.scala 31:69]
  wire [4:0] _T_370; // @[Mux.scala 31:69]
  wire [4:0] _T_371; // @[Mux.scala 31:69]
  wire [4:0] _T_372; // @[Mux.scala 31:69]
  wire [4:0] _T_373; // @[Mux.scala 31:69]
  wire [4:0] _T_374; // @[Mux.scala 31:69]
  wire [4:0] _T_375; // @[Mux.scala 31:69]
  wire [53:0] _GEN_39; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_376; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_378; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_40; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_379; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_380; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_381; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_41; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_382; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_42; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_384; // @[rawFloatFromFN.scala 59:15]
  wire  _T_385; // @[rawFloatFromFN.scala 62:34]
  wire  _T_387; // @[rawFloatFromFN.scala 63:62]
  wire  _T_391; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_394; // @[rawFloatFromFN.scala 70:48]
  wire [22:0] _T_396; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_398; // @[Cat.scala 30:58]
  wire [2:0] _T_400; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_43; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_402; // @[recFNFromFN.scala 48:79]
  wire [32:0] _T_407; // @[Cat.scala 30:58]
  wire  _T_411; // @[FPU.scala 265:42]
  wire [64:0] _T_422; // @[Cat.scala 30:58]
  wire  _T_425; // @[FPU.scala 197:56]
  wire [32:0] _T_434; // @[FPU.scala 473:45]
  wire [31:0] _T_435; // @[FPU.scala 473:60]
  wire [32:0] _T_436; // @[FPU.scala 473:19]
  wire [64:0] _T_442; // @[FPU.scala 340:25]
  wire  _T_445; // @[FPU.scala 197:56]
  wire [64:0] _T_446; // @[FPU.scala 341:10]
  wire [64:0] _T_448; // @[Cat.scala 30:58]
  reg [64:0] _T_456_data; // @[Reg.scala 11:16]
  reg [95:0] _RAND_6;
  reg [4:0] _T_456_exc; // @[Reg.scala 11:16]
  reg [31:0] _RAND_7;
  reg [4:0] IntToFP_state; // @[Register tracking IntToFP state]
  reg [31:0] _RAND_8;
  reg  IntToFP_cov [0:31]; // @[Coverage map for IntToFP]
  reg [31:0] _RAND_9;
  wire  IntToFP_cov_read_data; // @[Coverage map for IntToFP]
  wire [4:0] IntToFP_cov_read_addr; // @[Coverage map for IntToFP]
  wire  IntToFP_cov_write_data; // @[Coverage map for IntToFP]
  wire [4:0] IntToFP_cov_write_addr; // @[Coverage map for IntToFP]
  wire  IntToFP_cov_write_mask; // @[Coverage map for IntToFP]
  wire  IntToFP_cov_write_en; // @[Coverage map for IntToFP]
  reg [29:0] IntToFP_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_10;
  wire [1:0] in_bits_typ_shl;
  wire [4:0] in_bits_typ_pad;
  wire [2:0] in_bits_singleIn_shl;
  wire [4:0] in_bits_singleIn_pad;
  wire [3:0] in_valid_shl;
  wire [4:0] in_valid_pad;
  wire [4:0] in_bits_wflags_shl;
  wire [4:0] in_bits_wflags_pad;
  wire [4:0] IntToFP_xor1;
  wire [4:0] IntToFP_xor2;
  wire [4:0] IntToFP_xor0;
  wire [29:0] INToRecFN_sum;
  wire [29:0] INToRecFN_1_sum;
  wire  INToRecFN_metaAssert_wire;
  wire  INToRecFN_1_metaAssert_wire;
  wire  IntToFP_or0;
  reg  IntToFP_metaAssert;
  reg [31:0] _RAND_11;
  INToRecFN INToRecFN ( // @[FPU.scala 483:23]
    .io_signedIn(INToRecFN_io_signedIn),
    .io_in(INToRecFN_io_in),
    .io_roundingMode(INToRecFN_io_roundingMode),
    .io_out(INToRecFN_io_out),
    .io_exceptionFlags(INToRecFN_io_exceptionFlags),
    .io_covSum(INToRecFN_io_covSum),
    .metaAssert(INToRecFN_metaAssert)
  );
  INToRecFN_1 INToRecFN_1 ( // @[FPU.scala 483:23]
    .io_signedIn(INToRecFN_1_io_signedIn),
    .io_in(INToRecFN_1_io_in),
    .io_roundingMode(INToRecFN_1_io_roundingMode),
    .io_out(INToRecFN_1_io_out),
    .io_exceptionFlags(INToRecFN_1_io_exceptionFlags),
    .io_covSum(INToRecFN_1_io_covSum),
    .metaAssert(INToRecFN_1_metaAssert)
  );
  assign tag = ~in_bits_singleIn; // @[FPU.scala 462:13]
  assign _T_21 = tag ? 64'h0 : 64'hffffffff00000000; // @[package.scala 31:71]
  assign _T_22 = _T_21 | in_bits_in1; // @[FPU.scala 358:23]
  assign _T_26 = _T_22[62:52] == 11'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_27 = _T_22[51:0] == 52'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_32 = {{16'd0}, _T_22[31:16]}; // @[Bitwise.scala 103:31]
  assign _T_34 = {_T_22[15:0], 16'h0}; // @[Bitwise.scala 103:65]
  assign _T_36 = _T_34 & 32'hffff0000; // @[Bitwise.scala 103:75]
  assign _T_37 = _T_32 | _T_36; // @[Bitwise.scala 103:39]
  assign _GEN_24 = {{8'd0}, _T_37[31:8]}; // @[Bitwise.scala 103:31]
  assign _T_42 = _GEN_24 & 32'hff00ff; // @[Bitwise.scala 103:31]
  assign _T_44 = {_T_37[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_46 = _T_44 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  assign _T_47 = _T_42 | _T_46; // @[Bitwise.scala 103:39]
  assign _GEN_25 = {{4'd0}, _T_47[31:4]}; // @[Bitwise.scala 103:31]
  assign _T_52 = _GEN_25 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  assign _T_54 = {_T_47[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_56 = _T_54 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  assign _T_57 = _T_52 | _T_56; // @[Bitwise.scala 103:39]
  assign _GEN_26 = {{2'd0}, _T_57[31:2]}; // @[Bitwise.scala 103:31]
  assign _T_62 = _GEN_26 & 32'h33333333; // @[Bitwise.scala 103:31]
  assign _T_64 = {_T_57[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_66 = _T_64 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  assign _T_67 = _T_62 | _T_66; // @[Bitwise.scala 103:39]
  assign _GEN_27 = {{1'd0}, _T_67[31:1]}; // @[Bitwise.scala 103:31]
  assign _T_72 = _GEN_27 & 32'h55555555; // @[Bitwise.scala 103:31]
  assign _T_74 = {_T_67[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_76 = _T_74 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  assign _T_77 = _T_72 | _T_76; // @[Bitwise.scala 103:39]
  assign _T_83 = {{8'd0}, _T_22[47:40]}; // @[Bitwise.scala 103:31]
  assign _T_85 = {_T_22[39:32], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_87 = _T_85 & 16'hff00; // @[Bitwise.scala 103:75]
  assign _T_88 = _T_83 | _T_87; // @[Bitwise.scala 103:39]
  assign _GEN_28 = {{4'd0}, _T_88[15:4]}; // @[Bitwise.scala 103:31]
  assign _T_93 = _GEN_28 & 16'hf0f; // @[Bitwise.scala 103:31]
  assign _T_95 = {_T_88[11:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_97 = _T_95 & 16'hf0f0; // @[Bitwise.scala 103:75]
  assign _T_98 = _T_93 | _T_97; // @[Bitwise.scala 103:39]
  assign _GEN_29 = {{2'd0}, _T_98[15:2]}; // @[Bitwise.scala 103:31]
  assign _T_103 = _GEN_29 & 16'h3333; // @[Bitwise.scala 103:31]
  assign _T_105 = {_T_98[13:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_107 = _T_105 & 16'hcccc; // @[Bitwise.scala 103:75]
  assign _T_108 = _T_103 | _T_107; // @[Bitwise.scala 103:39]
  assign _GEN_30 = {{1'd0}, _T_108[15:1]}; // @[Bitwise.scala 103:31]
  assign _T_113 = _GEN_30 & 16'h5555; // @[Bitwise.scala 103:31]
  assign _T_115 = {_T_108[14:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_117 = _T_115 & 16'haaaa; // @[Bitwise.scala 103:75]
  assign _T_118 = _T_113 | _T_117; // @[Bitwise.scala 103:39]
  assign _T_130 = {_T_77,_T_118,_T_22[48],_T_22[49],_T_22[50],_T_22[51]}; // @[Cat.scala 30:58]
  assign _T_183 = _T_130[50] ? 6'h32 : 6'h33; // @[Mux.scala 31:69]
  assign _T_184 = _T_130[49] ? 6'h31 : _T_183; // @[Mux.scala 31:69]
  assign _T_185 = _T_130[48] ? 6'h30 : _T_184; // @[Mux.scala 31:69]
  assign _T_186 = _T_130[47] ? 6'h2f : _T_185; // @[Mux.scala 31:69]
  assign _T_187 = _T_130[46] ? 6'h2e : _T_186; // @[Mux.scala 31:69]
  assign _T_188 = _T_130[45] ? 6'h2d : _T_187; // @[Mux.scala 31:69]
  assign _T_189 = _T_130[44] ? 6'h2c : _T_188; // @[Mux.scala 31:69]
  assign _T_190 = _T_130[43] ? 6'h2b : _T_189; // @[Mux.scala 31:69]
  assign _T_191 = _T_130[42] ? 6'h2a : _T_190; // @[Mux.scala 31:69]
  assign _T_192 = _T_130[41] ? 6'h29 : _T_191; // @[Mux.scala 31:69]
  assign _T_193 = _T_130[40] ? 6'h28 : _T_192; // @[Mux.scala 31:69]
  assign _T_194 = _T_130[39] ? 6'h27 : _T_193; // @[Mux.scala 31:69]
  assign _T_195 = _T_130[38] ? 6'h26 : _T_194; // @[Mux.scala 31:69]
  assign _T_196 = _T_130[37] ? 6'h25 : _T_195; // @[Mux.scala 31:69]
  assign _T_197 = _T_130[36] ? 6'h24 : _T_196; // @[Mux.scala 31:69]
  assign _T_198 = _T_130[35] ? 6'h23 : _T_197; // @[Mux.scala 31:69]
  assign _T_199 = _T_130[34] ? 6'h22 : _T_198; // @[Mux.scala 31:69]
  assign _T_200 = _T_130[33] ? 6'h21 : _T_199; // @[Mux.scala 31:69]
  assign _T_201 = _T_130[32] ? 6'h20 : _T_200; // @[Mux.scala 31:69]
  assign _T_202 = _T_130[31] ? 6'h1f : _T_201; // @[Mux.scala 31:69]
  assign _T_203 = _T_130[30] ? 6'h1e : _T_202; // @[Mux.scala 31:69]
  assign _T_204 = _T_130[29] ? 6'h1d : _T_203; // @[Mux.scala 31:69]
  assign _T_205 = _T_130[28] ? 6'h1c : _T_204; // @[Mux.scala 31:69]
  assign _T_206 = _T_130[27] ? 6'h1b : _T_205; // @[Mux.scala 31:69]
  assign _T_207 = _T_130[26] ? 6'h1a : _T_206; // @[Mux.scala 31:69]
  assign _T_208 = _T_130[25] ? 6'h19 : _T_207; // @[Mux.scala 31:69]
  assign _T_209 = _T_130[24] ? 6'h18 : _T_208; // @[Mux.scala 31:69]
  assign _T_210 = _T_130[23] ? 6'h17 : _T_209; // @[Mux.scala 31:69]
  assign _T_211 = _T_130[22] ? 6'h16 : _T_210; // @[Mux.scala 31:69]
  assign _T_212 = _T_130[21] ? 6'h15 : _T_211; // @[Mux.scala 31:69]
  assign _T_213 = _T_130[20] ? 6'h14 : _T_212; // @[Mux.scala 31:69]
  assign _T_214 = _T_130[19] ? 6'h13 : _T_213; // @[Mux.scala 31:69]
  assign _T_215 = _T_130[18] ? 6'h12 : _T_214; // @[Mux.scala 31:69]
  assign _T_216 = _T_130[17] ? 6'h11 : _T_215; // @[Mux.scala 31:69]
  assign _T_217 = _T_130[16] ? 6'h10 : _T_216; // @[Mux.scala 31:69]
  assign _T_218 = _T_130[15] ? 6'hf : _T_217; // @[Mux.scala 31:69]
  assign _T_219 = _T_130[14] ? 6'he : _T_218; // @[Mux.scala 31:69]
  assign _T_220 = _T_130[13] ? 6'hd : _T_219; // @[Mux.scala 31:69]
  assign _T_221 = _T_130[12] ? 6'hc : _T_220; // @[Mux.scala 31:69]
  assign _T_222 = _T_130[11] ? 6'hb : _T_221; // @[Mux.scala 31:69]
  assign _T_223 = _T_130[10] ? 6'ha : _T_222; // @[Mux.scala 31:69]
  assign _T_224 = _T_130[9] ? 6'h9 : _T_223; // @[Mux.scala 31:69]
  assign _T_225 = _T_130[8] ? 6'h8 : _T_224; // @[Mux.scala 31:69]
  assign _T_226 = _T_130[7] ? 6'h7 : _T_225; // @[Mux.scala 31:69]
  assign _T_227 = _T_130[6] ? 6'h6 : _T_226; // @[Mux.scala 31:69]
  assign _T_228 = _T_130[5] ? 6'h5 : _T_227; // @[Mux.scala 31:69]
  assign _T_229 = _T_130[4] ? 6'h4 : _T_228; // @[Mux.scala 31:69]
  assign _T_230 = _T_130[3] ? 6'h3 : _T_229; // @[Mux.scala 31:69]
  assign _T_231 = _T_130[2] ? 6'h2 : _T_230; // @[Mux.scala 31:69]
  assign _T_232 = _T_130[1] ? 6'h1 : _T_231; // @[Mux.scala 31:69]
  assign _T_233 = _T_130[0] ? 6'h0 : _T_232; // @[Mux.scala 31:69]
  assign _GEN_31 = {{63'd0}, _T_22[51:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_234 = _GEN_31 << _T_233; // @[rawFloatFromFN.scala 54:36]
  assign _T_236 = {_T_234[50:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_32 = {{6'd0}, _T_233}; // @[rawFloatFromFN.scala 57:26]
  assign _T_237 = _GEN_32 ^ 12'hfff; // @[rawFloatFromFN.scala 57:26]
  assign _T_238 = _T_26 ? _T_237 : {{1'd0}, _T_22[62:52]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_239 = _T_26 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_33 = {{9'd0}, _T_239}; // @[rawFloatFromFN.scala 60:22]
  assign _T_240 = 11'h400 | _GEN_33; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_34 = {{1'd0}, _T_240}; // @[rawFloatFromFN.scala 59:15]
  assign _T_242 = _T_238 + _GEN_34; // @[rawFloatFromFN.scala 59:15]
  assign _T_243 = _T_26 & _T_27; // @[rawFloatFromFN.scala 62:34]
  assign _T_245 = _T_242[11:10] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_249 = _T_245 & ~_T_27; // @[rawFloatFromFN.scala 66:33]
  assign _T_252 = {1'b0,$signed(_T_242)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_254 = _T_26 ? _T_236 : _T_22[51:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_256 = {1'h0,~_T_243,_T_254}; // @[Cat.scala 30:58]
  assign _T_258 = _T_243 ? 3'h0 : _T_252[11:9]; // @[recFNFromFN.scala 48:16]
  assign _GEN_35 = {{2'd0}, _T_249}; // @[recFNFromFN.scala 48:79]
  assign _T_260 = _T_258 | _GEN_35; // @[recFNFromFN.scala 48:79]
  assign _T_265 = {_T_22[63],_T_260,_T_252[8:0],_T_256[51:0]}; // @[Cat.scala 30:58]
  assign _T_269 = _T_22[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_270 = _T_22[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_275 = {{8'd0}, _T_22[15:8]}; // @[Bitwise.scala 103:31]
  assign _T_277 = {_T_22[7:0], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_279 = _T_277 & 16'hff00; // @[Bitwise.scala 103:75]
  assign _T_280 = _T_275 | _T_279; // @[Bitwise.scala 103:39]
  assign _GEN_36 = {{4'd0}, _T_280[15:4]}; // @[Bitwise.scala 103:31]
  assign _T_285 = _GEN_36 & 16'hf0f; // @[Bitwise.scala 103:31]
  assign _T_287 = {_T_280[11:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_289 = _T_287 & 16'hf0f0; // @[Bitwise.scala 103:75]
  assign _T_290 = _T_285 | _T_289; // @[Bitwise.scala 103:39]
  assign _GEN_37 = {{2'd0}, _T_290[15:2]}; // @[Bitwise.scala 103:31]
  assign _T_295 = _GEN_37 & 16'h3333; // @[Bitwise.scala 103:31]
  assign _T_297 = {_T_290[13:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_299 = _T_297 & 16'hcccc; // @[Bitwise.scala 103:75]
  assign _T_300 = _T_295 | _T_299; // @[Bitwise.scala 103:39]
  assign _GEN_38 = {{1'd0}, _T_300[15:1]}; // @[Bitwise.scala 103:31]
  assign _T_305 = _GEN_38 & 16'h5555; // @[Bitwise.scala 103:31]
  assign _T_307 = {_T_300[14:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_309 = _T_307 & 16'haaaa; // @[Bitwise.scala 103:75]
  assign _T_310 = _T_305 | _T_309; // @[Bitwise.scala 103:39]
  assign _T_330 = {_T_310,_T_22[16],_T_22[17],_T_22[18],_T_22[19],_T_22[20],_T_22[21],_T_22[22]}; // @[Cat.scala 30:58]
  assign _T_354 = _T_330[21] ? 5'h15 : 5'h16; // @[Mux.scala 31:69]
  assign _T_355 = _T_330[20] ? 5'h14 : _T_354; // @[Mux.scala 31:69]
  assign _T_356 = _T_330[19] ? 5'h13 : _T_355; // @[Mux.scala 31:69]
  assign _T_357 = _T_330[18] ? 5'h12 : _T_356; // @[Mux.scala 31:69]
  assign _T_358 = _T_330[17] ? 5'h11 : _T_357; // @[Mux.scala 31:69]
  assign _T_359 = _T_330[16] ? 5'h10 : _T_358; // @[Mux.scala 31:69]
  assign _T_360 = _T_330[15] ? 5'hf : _T_359; // @[Mux.scala 31:69]
  assign _T_361 = _T_330[14] ? 5'he : _T_360; // @[Mux.scala 31:69]
  assign _T_362 = _T_330[13] ? 5'hd : _T_361; // @[Mux.scala 31:69]
  assign _T_363 = _T_330[12] ? 5'hc : _T_362; // @[Mux.scala 31:69]
  assign _T_364 = _T_330[11] ? 5'hb : _T_363; // @[Mux.scala 31:69]
  assign _T_365 = _T_330[10] ? 5'ha : _T_364; // @[Mux.scala 31:69]
  assign _T_366 = _T_330[9] ? 5'h9 : _T_365; // @[Mux.scala 31:69]
  assign _T_367 = _T_330[8] ? 5'h8 : _T_366; // @[Mux.scala 31:69]
  assign _T_368 = _T_330[7] ? 5'h7 : _T_367; // @[Mux.scala 31:69]
  assign _T_369 = _T_330[6] ? 5'h6 : _T_368; // @[Mux.scala 31:69]
  assign _T_370 = _T_330[5] ? 5'h5 : _T_369; // @[Mux.scala 31:69]
  assign _T_371 = _T_330[4] ? 5'h4 : _T_370; // @[Mux.scala 31:69]
  assign _T_372 = _T_330[3] ? 5'h3 : _T_371; // @[Mux.scala 31:69]
  assign _T_373 = _T_330[2] ? 5'h2 : _T_372; // @[Mux.scala 31:69]
  assign _T_374 = _T_330[1] ? 5'h1 : _T_373; // @[Mux.scala 31:69]
  assign _T_375 = _T_330[0] ? 5'h0 : _T_374; // @[Mux.scala 31:69]
  assign _GEN_39 = {{31'd0}, _T_22[22:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_376 = _GEN_39 << _T_375; // @[rawFloatFromFN.scala 54:36]
  assign _T_378 = {_T_376[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_40 = {{4'd0}, _T_375}; // @[rawFloatFromFN.scala 57:26]
  assign _T_379 = _GEN_40 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  assign _T_380 = _T_269 ? _T_379 : {{1'd0}, _T_22[30:23]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_381 = _T_269 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_41 = {{6'd0}, _T_381}; // @[rawFloatFromFN.scala 60:22]
  assign _T_382 = 8'h80 | _GEN_41; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_42 = {{1'd0}, _T_382}; // @[rawFloatFromFN.scala 59:15]
  assign _T_384 = _T_380 + _GEN_42; // @[rawFloatFromFN.scala 59:15]
  assign _T_385 = _T_269 & _T_270; // @[rawFloatFromFN.scala 62:34]
  assign _T_387 = _T_384[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_391 = _T_387 & ~_T_270; // @[rawFloatFromFN.scala 66:33]
  assign _T_394 = {1'b0,$signed(_T_384)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_396 = _T_269 ? _T_378 : _T_22[22:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_398 = {1'h0,~_T_385,_T_396}; // @[Cat.scala 30:58]
  assign _T_400 = _T_385 ? 3'h0 : _T_394[8:6]; // @[recFNFromFN.scala 48:16]
  assign _GEN_43 = {{2'd0}, _T_391}; // @[recFNFromFN.scala 48:79]
  assign _T_402 = _T_400 | _GEN_43; // @[recFNFromFN.scala 48:79]
  assign _T_407 = {_T_22[31],_T_402,_T_394[5:0],_T_398[22:0]}; // @[Cat.scala 30:58]
  assign _T_411 = ~_T_265[51:32] == 20'h0; // @[FPU.scala 265:42]
  assign _T_422 = {_T_265[64:61],_T_411,_T_265[59:53],_T_407[31],_T_265[51:32],_T_407[32],_T_407[30:0]}; // @[Cat.scala 30:58]
  assign _T_425 = ~_T_265[63:61] == 3'h0; // @[FPU.scala 197:56]
  assign _T_434 = {1'b0,$signed(in_bits_in1[31:0])}; // @[FPU.scala 473:45]
  assign _T_435 = in_bits_in1[31:0]; // @[FPU.scala 473:60]
  assign _T_436 = in_bits_typ[0] ? $signed(_T_434) : $signed({{1{_T_435[31]}},_T_435}); // @[FPU.scala 473:19]
  assign _T_442 = INToRecFN_1_io_out & 65'h1efefffffffffffff; // @[FPU.scala 340:25]
  assign _T_445 = ~INToRecFN_1_io_out[63:61] == 3'h0; // @[FPU.scala 197:56]
  assign _T_446 = _T_445 ? _T_442 : INToRecFN_1_io_out; // @[FPU.scala 341:10]
  assign _T_448 = {_T_446[64:33],INToRecFN_io_out}; // @[Cat.scala 30:58]
  assign io_out_bits_data = _T_456_data; // @[FPU.scala 497:10]
  assign io_out_bits_exc = _T_456_exc; // @[FPU.scala 497:10]
  assign INToRecFN_io_signedIn = ~in_bits_typ[0]; // @[FPU.scala 484:23]
  assign INToRecFN_io_in = in_bits_typ[1] ? $signed(in_bits_in1) : $signed({{31{_T_436[32]}},_T_436}); // @[FPU.scala 485:17]
  assign INToRecFN_io_roundingMode = in_bits_rm; // @[FPU.scala 486:27]
  assign INToRecFN_1_io_signedIn = ~in_bits_typ[0]; // @[FPU.scala 484:23]
  assign INToRecFN_1_io_in = in_bits_typ[1] ? $signed(in_bits_in1) : $signed({{31{_T_436[32]}},_T_436}); // @[FPU.scala 485:17]
  assign INToRecFN_1_io_roundingMode = in_bits_rm; // @[FPU.scala 486:27]
  assign IntToFP_cov_read_addr = IntToFP_state;
  assign IntToFP_cov_read_data = IntToFP_cov[IntToFP_cov_read_addr]; // @[Coverage map for IntToFP]
  assign IntToFP_cov_write_data = 1'h1;
  assign IntToFP_cov_write_addr = IntToFP_state;
  assign IntToFP_cov_write_mask = 1'h1;
  assign IntToFP_cov_write_en = 1'h1;
  assign in_bits_typ_shl = in_bits_typ;
  assign in_bits_typ_pad = {3'h0,in_bits_typ_shl};
  assign in_bits_singleIn_shl = {in_bits_singleIn, 2'h0};
  assign in_bits_singleIn_pad = {2'h0,in_bits_singleIn_shl};
  assign in_valid_shl = {in_valid, 3'h0};
  assign in_valid_pad = {1'h0,in_valid_shl};
  assign in_bits_wflags_shl = {in_bits_wflags, 4'h0};
  assign in_bits_wflags_pad = in_bits_wflags_shl;
  assign IntToFP_xor1 = in_bits_typ_pad ^ in_bits_singleIn_pad;
  assign IntToFP_xor2 = in_valid_pad ^ in_bits_wflags_pad;
  assign IntToFP_xor0 = IntToFP_xor1 ^ IntToFP_xor2;
  assign INToRecFN_sum = IntToFP_covSum + INToRecFN_io_covSum;
  assign INToRecFN_1_sum = INToRecFN_sum + INToRecFN_1_io_covSum;
  assign io_covSum = INToRecFN_1_sum;
  assign INToRecFN_metaAssert_wire = INToRecFN_metaAssert;
  assign INToRecFN_1_metaAssert_wire = INToRecFN_1_metaAssert;
  assign IntToFP_or0 = INToRecFN_metaAssert_wire | INToRecFN_1_metaAssert_wire;
  assign metaAssert = IntToFP_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_bits_singleIn = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_bits_wflags = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_bits_rm = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  in_bits_typ = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {2{`RANDOM}};
  in_bits_in1 = _RAND_5[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {3{`RANDOM}};
  _T_456_data = _RAND_6[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_456_exc = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  IntToFP_state = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    IntToFP_cov[initvar] = _RAND_9[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  IntToFP_covSum = _RAND_10[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  IntToFP_metaAssert = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      in_valid <= 1'h0;
    end else if (reset) begin
      in_valid <= 1'h0;
    end else begin
      in_valid <= io_in_valid;
    end
    if (metaReset) begin
      in_bits_singleIn <= 1'h0;
    end else if (io_in_valid) begin
      in_bits_singleIn <= io_in_bits_singleIn;
    end
    if (metaReset) begin
      in_bits_wflags <= 1'h0;
    end else if (io_in_valid) begin
      in_bits_wflags <= io_in_bits_wflags;
    end
    if (metaReset) begin
      in_bits_rm <= 3'h0;
    end else if (io_in_valid) begin
      in_bits_rm <= io_in_bits_rm;
    end
    if (metaReset) begin
      in_bits_typ <= 2'h0;
    end else if (io_in_valid) begin
      in_bits_typ <= io_in_bits_typ;
    end
    if (metaReset) begin
      in_bits_in1 <= 64'h0;
    end else if (io_in_valid) begin
      in_bits_in1 <= io_in_bits_in1;
    end
    if (metaReset) begin
      _T_456_data <= 65'h0;
    end else if (in_valid) begin
      if (in_bits_wflags) begin
        if (tag) begin
          if (_T_445) begin
            _T_456_data <= _T_442;
          end else begin
            _T_456_data <= INToRecFN_1_io_out;
          end
        end else begin
          _T_456_data <= _T_448;
        end
      end else if (_T_425) begin
        _T_456_data <= _T_422;
      end else begin
        _T_456_data <= _T_265;
      end
    end
    if (metaReset) begin
      _T_456_exc <= 5'h0;
    end else if (in_valid) begin
      if (in_bits_wflags) begin
        if (tag) begin
          _T_456_exc <= INToRecFN_1_io_exceptionFlags;
        end else begin
          _T_456_exc <= INToRecFN_io_exceptionFlags;
        end
      end else begin
        _T_456_exc <= 5'h0;
      end
    end
    IntToFP_state <= IntToFP_xor0;
    if (!(IntToFP_cov_read_data)) begin
      IntToFP_covSum <= IntToFP_covSum + 1'h1;
    end
    if (metaReset) begin
      IntToFP_metaAssert <= 1'h0;
    end else begin
      IntToFP_metaAssert <= IntToFP_metaAssert | IntToFP_or0;
    end
  end
  always @(posedge clock) begin
    if(IntToFP_cov_write_en & IntToFP_cov_write_mask) begin
      IntToFP_cov[IntToFP_cov_write_addr] <= IntToFP_cov_write_data; // @[Coverage map for IntToFP]
    end
  end
endmodule
module FPToFP(
  input         clock,
  input         reset,
  input         io_in_valid,
  input         io_in_bits_ren2,
  input         io_in_bits_singleOut,
  input         io_in_bits_wflags,
  input  [2:0]  io_in_bits_rm,
  input  [64:0] io_in_bits_in1,
  input  [64:0] io_in_bits_in2,
  output [64:0] io_out_bits_data,
  output [4:0]  io_out_bits_exc,
  input         io_lt,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [64:0] RecFNToRecFN_io_in; // @[FPU.scala 546:30]
  wire [2:0] RecFNToRecFN_io_roundingMode; // @[FPU.scala 546:30]
  wire [32:0] RecFNToRecFN_io_out; // @[FPU.scala 546:30]
  wire [4:0] RecFNToRecFN_io_exceptionFlags; // @[FPU.scala 546:30]
  wire [29:0] RecFNToRecFN_io_covSum; // @[FPU.scala 546:30]
  wire  RecFNToRecFN_metaAssert; // @[FPU.scala 546:30]
  reg  in_valid; // @[Valid.scala 48:22]
  reg [31:0] _RAND_0;
  reg  in_bits_ren2; // @[Reg.scala 11:16]
  reg [31:0] _RAND_1;
  reg  in_bits_singleOut; // @[Reg.scala 11:16]
  reg [31:0] _RAND_2;
  reg  in_bits_wflags; // @[Reg.scala 11:16]
  reg [31:0] _RAND_3;
  reg [2:0] in_bits_rm; // @[Reg.scala 11:16]
  reg [31:0] _RAND_4;
  reg [64:0] in_bits_in1; // @[Reg.scala 11:16]
  reg [95:0] _RAND_5;
  reg [64:0] in_bits_in2; // @[Reg.scala 11:16]
  reg [95:0] _RAND_6;
  wire [64:0] _T_20; // @[FPU.scala 509:48]
  wire [64:0] _T_23; // @[FPU.scala 509:66]
  wire [64:0] signNum; // @[FPU.scala 509:20]
  wire [64:0] fsgnj; // @[Cat.scala 30:58]
  wire  _T_29; // @[FPU.scala 197:56]
  wire  _T_32; // @[FPU.scala 197:56]
  wire  _T_38; // @[FPU.scala 198:34]
  wire  _T_44; // @[FPU.scala 198:34]
  wire  _T_45; // @[FPU.scala 519:49]
  wire  _T_46; // @[FPU.scala 520:27]
  wire  _T_48; // @[FPU.scala 521:41]
  wire  _T_50; // @[FPU.scala 521:51]
  wire  _T_51; // @[FPU.scala 521:24]
  wire [4:0] _T_52; // @[FPU.scala 522:31]
  wire [64:0] _T_53; // @[FPU.scala 523:53]
  wire [64:0] _T_54; // @[FPU.scala 523:25]
  wire [64:0] _GEN_23; // @[FPU.scala 516:25]
  wire  outTag; // @[FPU.scala 527:16]
  wire  _T_80; // @[FPU.scala 535:24]
  wire [64:0] _T_84; // @[FPU.scala 538:24]
  wire [64:0] fsgnjMux_data; // @[FPU.scala 535:42]
  wire [75:0] _T_61; // @[FPU.scala 225:28]
  wire [11:0] _T_65; // @[FPU.scala 228:31]
  wire [11:0] _T_68; // @[FPU.scala 228:48]
  wire  _T_69; // @[FPU.scala 229:19]
  wire  _T_70; // @[FPU.scala 229:36]
  wire  _T_71; // @[FPU.scala 229:25]
  wire [8:0] _T_73; // @[Cat.scala 30:58]
  wire [8:0] _T_75; // @[FPU.scala 229:10]
  wire [64:0] _T_78; // @[Cat.scala 30:58]
  wire [4:0] _T_91; // @[FPU.scala 540:51]
  wire [64:0] _T_97; // @[Cat.scala 30:58]
  reg [64:0] _T_101_data; // @[Reg.scala 11:16]
  reg [95:0] _RAND_7;
  reg [4:0] _T_101_exc; // @[Reg.scala 11:16]
  reg [31:0] _RAND_8;
  reg [6:0] FPToFP_state; // @[Register tracking FPToFP state]
  reg [31:0] _RAND_9;
  reg  FPToFP_cov [0:127]; // @[Coverage map for FPToFP]
  reg [31:0] _RAND_10;
  wire  FPToFP_cov_read_data; // @[Coverage map for FPToFP]
  wire [6:0] FPToFP_cov_read_addr; // @[Coverage map for FPToFP]
  wire  FPToFP_cov_write_data; // @[Coverage map for FPToFP]
  wire [6:0] FPToFP_cov_write_addr; // @[Coverage map for FPToFP]
  wire  FPToFP_cov_write_mask; // @[Coverage map for FPToFP]
  wire  FPToFP_cov_write_en; // @[Coverage map for FPToFP]
  reg [29:0] FPToFP_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_11;
  wire  in_bits_singleOut_shl;
  wire [6:0] in_bits_singleOut_pad;
  wire [1:0] in_valid_shl;
  wire [6:0] in_valid_pad;
  wire [2:0] in_bits_ren2_shl;
  wire [6:0] in_bits_ren2_pad;
  wire [3:0] in_bits_wflags_shl;
  wire [6:0] in_bits_wflags_pad;
  wire [6:0] in_bits_rm_shl;
  wire [6:0] in_bits_rm_pad;
  wire [6:0] FPToFP_xor1;
  wire [6:0] FPToFP_xor6;
  wire [6:0] FPToFP_xor2;
  wire [6:0] FPToFP_xor0;
  wire [29:0] RecFNToRecFN_sum;
  wire  RecFNToRecFN_metaAssert_wire;
  reg  FPToFP_metaAssert;
  reg [31:0] _RAND_12;
  RecFNToRecFN RecFNToRecFN ( // @[FPU.scala 546:30]
    .io_in(RecFNToRecFN_io_in),
    .io_roundingMode(RecFNToRecFN_io_roundingMode),
    .io_out(RecFNToRecFN_io_out),
    .io_exceptionFlags(RecFNToRecFN_io_exceptionFlags),
    .io_covSum(RecFNToRecFN_io_covSum),
    .metaAssert(RecFNToRecFN_metaAssert)
  );
  assign _T_20 = in_bits_in1 ^ in_bits_in2; // @[FPU.scala 509:48]
  assign _T_23 = in_bits_rm[0] ? ~in_bits_in2 : in_bits_in2; // @[FPU.scala 509:66]
  assign signNum = in_bits_rm[1] ? _T_20 : _T_23; // @[FPU.scala 509:20]
  assign fsgnj = {signNum[64],in_bits_in1[63:0]}; // @[Cat.scala 30:58]
  assign _T_29 = ~in_bits_in1[63:61] == 3'h0; // @[FPU.scala 197:56]
  assign _T_32 = ~in_bits_in2[63:61] == 3'h0; // @[FPU.scala 197:56]
  assign _T_38 = _T_29 & ~in_bits_in1[51]; // @[FPU.scala 198:34]
  assign _T_44 = _T_32 & ~in_bits_in2[51]; // @[FPU.scala 198:34]
  assign _T_45 = _T_38 | _T_44; // @[FPU.scala 519:49]
  assign _T_46 = _T_29 & _T_32; // @[FPU.scala 520:27]
  assign _T_48 = in_bits_rm[0] != io_lt; // @[FPU.scala 521:41]
  assign _T_50 = _T_48 & ~_T_29; // @[FPU.scala 521:51]
  assign _T_51 = _T_32 | _T_50; // @[FPU.scala 521:24]
  assign _T_52 = {_T_45, 4'h0}; // @[FPU.scala 522:31]
  assign _T_53 = _T_51 ? in_bits_in1 : in_bits_in2; // @[FPU.scala 523:53]
  assign _T_54 = _T_46 ? 65'he008000000000000 : _T_53; // @[FPU.scala 523:25]
  assign _GEN_23 = in_bits_wflags ? _T_54 : fsgnj; // @[FPU.scala 516:25]
  assign outTag = ~in_bits_singleOut; // @[FPU.scala 527:16]
  assign _T_80 = in_bits_wflags & ~in_bits_ren2; // @[FPU.scala 535:24]
  assign _T_84 = _T_29 ? 65'he008000000000000 : in_bits_in1; // @[FPU.scala 538:24]
  assign fsgnjMux_data = _T_80 ? _T_84 : _GEN_23; // @[FPU.scala 535:42]
  assign _T_61 = {fsgnjMux_data[51:0], 24'h0}; // @[FPU.scala 225:28]
  assign _T_65 = fsgnjMux_data[63:52] + 12'h100; // @[FPU.scala 228:31]
  assign _T_68 = _T_65 - 12'h800; // @[FPU.scala 228:48]
  assign _T_69 = fsgnjMux_data[63:61] == 3'h0; // @[FPU.scala 229:19]
  assign _T_70 = fsgnjMux_data[63:61] >= 3'h6; // @[FPU.scala 229:36]
  assign _T_71 = _T_69 | _T_70; // @[FPU.scala 229:25]
  assign _T_73 = {fsgnjMux_data[63:61],_T_68[5:0]}; // @[Cat.scala 30:58]
  assign _T_75 = _T_71 ? _T_73 : _T_68[8:0]; // @[FPU.scala 229:10]
  assign _T_78 = {fsgnjMux_data[64:33],fsgnjMux_data[64],_T_75,_T_61[75:53]}; // @[Cat.scala 30:58]
  assign _T_91 = {_T_38, 4'h0}; // @[FPU.scala 540:51]
  assign _T_97 = {fsgnjMux_data[64:33],RecFNToRecFN_io_out}; // @[Cat.scala 30:58]
  assign io_out_bits_data = _T_101_data; // @[FPU.scala 557:10]
  assign io_out_bits_exc = _T_101_exc; // @[FPU.scala 557:10]
  assign RecFNToRecFN_io_in = in_bits_in1; // @[FPU.scala 547:24]
  assign RecFNToRecFN_io_roundingMode = in_bits_rm; // @[FPU.scala 548:34]
  assign FPToFP_cov_read_addr = FPToFP_state;
  assign FPToFP_cov_read_data = FPToFP_cov[FPToFP_cov_read_addr]; // @[Coverage map for FPToFP]
  assign FPToFP_cov_write_data = 1'h1;
  assign FPToFP_cov_write_addr = FPToFP_state;
  assign FPToFP_cov_write_mask = 1'h1;
  assign FPToFP_cov_write_en = 1'h1;
  assign in_bits_singleOut_shl = in_bits_singleOut;
  assign in_bits_singleOut_pad = {6'h0,in_bits_singleOut_shl};
  assign in_valid_shl = {in_valid, 1'h0};
  assign in_valid_pad = {5'h0,in_valid_shl};
  assign in_bits_ren2_shl = {in_bits_ren2, 2'h0};
  assign in_bits_ren2_pad = {4'h0,in_bits_ren2_shl};
  assign in_bits_wflags_shl = {in_bits_wflags, 3'h0};
  assign in_bits_wflags_pad = {3'h0,in_bits_wflags_shl};
  assign in_bits_rm_shl = {in_bits_rm, 4'h0};
  assign in_bits_rm_pad = in_bits_rm_shl;
  assign FPToFP_xor1 = in_bits_singleOut_pad ^ in_valid_pad;
  assign FPToFP_xor6 = in_bits_wflags_pad ^ in_bits_rm_pad;
  assign FPToFP_xor2 = in_bits_ren2_pad ^ FPToFP_xor6;
  assign FPToFP_xor0 = FPToFP_xor1 ^ FPToFP_xor2;
  assign RecFNToRecFN_sum = FPToFP_covSum + RecFNToRecFN_io_covSum;
  assign io_covSum = RecFNToRecFN_sum;
  assign RecFNToRecFN_metaAssert_wire = RecFNToRecFN_metaAssert;
  assign metaAssert = FPToFP_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_bits_ren2 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_bits_singleOut = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_bits_wflags = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  in_bits_rm = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {3{`RANDOM}};
  in_bits_in1 = _RAND_5[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {3{`RANDOM}};
  in_bits_in2 = _RAND_6[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {3{`RANDOM}};
  _T_101_data = _RAND_7[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_101_exc = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  FPToFP_state = _RAND_9[6:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    FPToFP_cov[initvar] = _RAND_10[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  FPToFP_covSum = _RAND_11[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  FPToFP_metaAssert = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      in_valid <= 1'h0;
    end else if (reset) begin
      in_valid <= 1'h0;
    end else begin
      in_valid <= io_in_valid;
    end
    if (metaReset) begin
      in_bits_ren2 <= 1'h0;
    end else if (io_in_valid) begin
      in_bits_ren2 <= io_in_bits_ren2;
    end
    if (metaReset) begin
      in_bits_singleOut <= 1'h0;
    end else if (io_in_valid) begin
      in_bits_singleOut <= io_in_bits_singleOut;
    end
    if (metaReset) begin
      in_bits_wflags <= 1'h0;
    end else if (io_in_valid) begin
      in_bits_wflags <= io_in_bits_wflags;
    end
    if (metaReset) begin
      in_bits_rm <= 3'h0;
    end else if (io_in_valid) begin
      in_bits_rm <= io_in_bits_rm;
    end
    if (metaReset) begin
      in_bits_in1 <= 65'h0;
    end else if (io_in_valid) begin
      in_bits_in1 <= io_in_bits_in1;
    end
    if (metaReset) begin
      in_bits_in2 <= 65'h0;
    end else if (io_in_valid) begin
      in_bits_in2 <= io_in_bits_in2;
    end
    if (metaReset) begin
      _T_101_data <= 65'h0;
    end else if (in_valid) begin
      if (_T_80) begin
        if (~outTag) begin
          _T_101_data <= _T_97;
        end else if (~outTag) begin
          _T_101_data <= _T_78;
        end else if (_T_80) begin
          if (_T_29) begin
            _T_101_data <= 65'he008000000000000;
          end else begin
            _T_101_data <= in_bits_in1;
          end
        end else if (in_bits_wflags) begin
          if (_T_46) begin
            _T_101_data <= 65'he008000000000000;
          end else if (_T_51) begin
            _T_101_data <= in_bits_in1;
          end else begin
            _T_101_data <= in_bits_in2;
          end
        end else begin
          _T_101_data <= fsgnj;
        end
      end else if (~outTag) begin
        _T_101_data <= _T_78;
      end else if (_T_80) begin
        if (_T_29) begin
          _T_101_data <= 65'he008000000000000;
        end else begin
          _T_101_data <= in_bits_in1;
        end
      end else if (in_bits_wflags) begin
        if (_T_46) begin
          _T_101_data <= 65'he008000000000000;
        end else if (_T_51) begin
          _T_101_data <= in_bits_in1;
        end else begin
          _T_101_data <= in_bits_in2;
        end
      end else begin
        _T_101_data <= fsgnj;
      end
    end
    if (metaReset) begin
      _T_101_exc <= 5'h0;
    end else if (in_valid) begin
      if (_T_80) begin
        if (~outTag) begin
          _T_101_exc <= RecFNToRecFN_io_exceptionFlags;
        end else if (_T_80) begin
          _T_101_exc <= _T_91;
        end else if (in_bits_wflags) begin
          _T_101_exc <= _T_52;
        end else begin
          _T_101_exc <= 5'h0;
        end
      end else if (_T_80) begin
        _T_101_exc <= _T_91;
      end else if (in_bits_wflags) begin
        _T_101_exc <= _T_52;
      end else begin
        _T_101_exc <= 5'h0;
      end
    end
    FPToFP_state <= FPToFP_xor0;
    if (!(FPToFP_cov_read_data)) begin
      FPToFP_covSum <= FPToFP_covSum + 1'h1;
    end
    if (metaReset) begin
      FPToFP_metaAssert <= 1'h0;
    end else begin
      FPToFP_metaAssert <= FPToFP_metaAssert | RecFNToRecFN_metaAssert_wire;
    end
  end
  always @(posedge clock) begin
    if(FPToFP_cov_write_en & FPToFP_cov_write_mask) begin
      FPToFP_cov[FPToFP_cov_write_addr] <= FPToFP_cov_write_data; // @[Coverage map for FPToFP]
    end
  end
endmodule
module FPUFMAPipe_1(
  input         clock,
  input         reset,
  input         io_in_valid,
  input         io_in_bits_ren3,
  input         io_in_bits_swap23,
  input  [2:0]  io_in_bits_rm,
  input  [1:0]  io_in_bits_fmaCmd,
  input  [64:0] io_in_bits_in1,
  input  [64:0] io_in_bits_in2,
  input  [64:0] io_in_bits_in3,
  output [64:0] io_out_bits_data,
  output [4:0]  io_out_bits_exc,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         fma_halt
);
  wire  fma_clock; // @[FPU.scala 644:19]
  wire  fma_reset; // @[FPU.scala 644:19]
  wire  fma_io_validin; // @[FPU.scala 644:19]
  wire [1:0] fma_io_op; // @[FPU.scala 644:19]
  wire [64:0] fma_io_a; // @[FPU.scala 644:19]
  wire [64:0] fma_io_b; // @[FPU.scala 644:19]
  wire [64:0] fma_io_c; // @[FPU.scala 644:19]
  wire [2:0] fma_io_roundingMode; // @[FPU.scala 644:19]
  wire [64:0] fma_io_out; // @[FPU.scala 644:19]
  wire [4:0] fma_io_exceptionFlags; // @[FPU.scala 644:19]
  wire  fma_io_validout; // @[FPU.scala 644:19]
  wire [29:0] fma_io_covSum; // @[FPU.scala 644:19]
  wire  fma_metaAssert; // @[FPU.scala 644:19]
  wire  fma_metaReset; // @[FPU.scala 644:19]
  reg  valid; // @[FPU.scala 632:18]
  reg [31:0] _RAND_0;
  reg [2:0] in_rm; // @[FPU.scala 633:15]
  reg [31:0] _RAND_1;
  reg [1:0] in_fmaCmd; // @[FPU.scala 633:15]
  reg [31:0] _RAND_2;
  reg [64:0] in_in1; // @[FPU.scala 633:15]
  reg [95:0] _RAND_3;
  reg [64:0] in_in2; // @[FPU.scala 633:15]
  reg [95:0] _RAND_4;
  reg [64:0] in_in3; // @[FPU.scala 633:15]
  reg [95:0] _RAND_5;
  wire [64:0] _T_13; // @[FPU.scala 636:32]
  wire [64:0] _T_15; // @[FPU.scala 636:50]
  wire  _T_16; // @[FPU.scala 641:21]
  wire [64:0] _T_20; // @[FPU.scala 340:25]
  wire  _T_23; // @[FPU.scala 197:56]
  reg [64:0] _T_28_data; // @[Reg.scala 11:16]
  reg [95:0] _RAND_6;
  reg [4:0] _T_28_exc; // @[Reg.scala 11:16]
  reg [31:0] _RAND_7;
  wire [4:0] res_exc; // @[FPU.scala 653:17 FPU.scala 655:11]
  wire [29:0] FPUFMAPipe_1_covSum;
  wire [29:0] fma_sum;
  wire  fma_metaAssert_wire;
  reg  FPUFMAPipe_1_metaAssert;
  reg [31:0] _RAND_8;
  MulAddRecFNPipe_1 fma ( // @[FPU.scala 644:19]
    .clock(fma_clock),
    .reset(fma_reset),
    .io_validin(fma_io_validin),
    .io_op(fma_io_op),
    .io_a(fma_io_a),
    .io_b(fma_io_b),
    .io_c(fma_io_c),
    .io_roundingMode(fma_io_roundingMode),
    .io_out(fma_io_out),
    .io_exceptionFlags(fma_io_exceptionFlags),
    .io_validout(fma_io_validout),
    .io_covSum(fma_io_covSum),
    .metaAssert(fma_metaAssert),
    .metaReset(fma_metaReset)
  );
  assign _T_13 = io_in_bits_in1 ^ io_in_bits_in2; // @[FPU.scala 636:32]
  assign _T_15 = _T_13 & 65'h10000000000000000; // @[FPU.scala 636:50]
  assign _T_16 = io_in_bits_ren3 | io_in_bits_swap23; // @[FPU.scala 641:21]
  assign _T_20 = fma_io_out & 65'h1efefffffffffffff; // @[FPU.scala 340:25]
  assign _T_23 = ~fma_io_out[63:61] == 3'h0; // @[FPU.scala 197:56]
  assign res_exc = fma_io_exceptionFlags; // @[FPU.scala 653:17 FPU.scala 655:11]
  assign io_out_bits_data = _T_28_data; // @[FPU.scala 657:10]
  assign io_out_bits_exc = _T_28_exc; // @[FPU.scala 657:10]
  assign fma_clock = clock;
  assign fma_reset = reset;
  assign fma_io_validin = valid; // @[FPU.scala 645:18]
  assign fma_io_op = in_fmaCmd; // @[FPU.scala 646:13]
  assign fma_io_a = in_in1; // @[FPU.scala 649:12]
  assign fma_io_b = in_in2; // @[FPU.scala 650:12]
  assign fma_io_c = in_in3; // @[FPU.scala 651:12]
  assign fma_io_roundingMode = in_rm; // @[FPU.scala 647:23]
  assign FPUFMAPipe_1_covSum = 30'h0;
  assign fma_sum = FPUFMAPipe_1_covSum + fma_io_covSum;
  assign io_covSum = fma_sum;
  assign fma_metaAssert_wire = fma_metaAssert;
  assign metaAssert = FPUFMAPipe_1_metaAssert;
  assign fma_metaReset = metaReset | fma_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_rm = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_fmaCmd = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {3{`RANDOM}};
  in_in1 = _RAND_3[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {3{`RANDOM}};
  in_in2 = _RAND_4[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {3{`RANDOM}};
  in_in3 = _RAND_5[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {3{`RANDOM}};
  _T_28_data = _RAND_6[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_28_exc = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  FPUFMAPipe_1_metaAssert = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      valid <= 1'h0;
    end else begin
      valid <= io_in_valid;
    end
    if (metaReset) begin
      in_rm <= 3'h0;
    end else if (io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if (metaReset) begin
      in_fmaCmd <= 2'h0;
    end else if (io_in_valid) begin
      in_fmaCmd <= io_in_bits_fmaCmd;
    end
    if (metaReset) begin
      in_in1 <= 65'h0;
    end else if (io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if (metaReset) begin
      in_in2 <= 65'h0;
    end else if (io_in_valid) begin
      if (io_in_bits_swap23) begin
        in_in2 <= 65'h8000000000000000;
      end else begin
        in_in2 <= io_in_bits_in2;
      end
    end
    if (metaReset) begin
      in_in3 <= 65'h0;
    end else if (io_in_valid) begin
      if (~_T_16) begin
        in_in3 <= _T_15;
      end else begin
        in_in3 <= io_in_bits_in3;
      end
    end
    if (metaReset) begin
      _T_28_data <= 65'h0;
    end else if (fma_io_validout) begin
      if (_T_23) begin
        _T_28_data <= _T_20;
      end else begin
        _T_28_data <= fma_io_out;
      end
    end
    if (metaReset) begin
      _T_28_exc <= 5'h0;
    end else if (fma_io_validout) begin
      _T_28_exc <= res_exc;
    end
    if (metaReset) begin
      FPUFMAPipe_1_metaAssert <= 1'h0;
    end else begin
      FPUFMAPipe_1_metaAssert <= FPUFMAPipe_1_metaAssert | fma_metaAssert_wire;
    end
  end
endmodule
module DivSqrtRecFN_small(
  input         clock,
  input         reset,
  output        io_inReady,
  input         io_inValid,
  input         io_sqrtOp,
  input  [32:0] io_a,
  input  [32:0] io_b,
  input  [2:0]  io_roundingMode,
  output        io_outValid_div,
  output        io_outValid_sqrt,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         divSqrtRecFNToRaw_halt
);
  wire  divSqrtRecFNToRaw_clock; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_reset; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_io_inReady; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_io_inValid; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_io_sqrtOp; // @[DivSqrtRecFN_small.scala 267:15]
  wire [32:0] divSqrtRecFNToRaw_io_a; // @[DivSqrtRecFN_small.scala 267:15]
  wire [32:0] divSqrtRecFNToRaw_io_b; // @[DivSqrtRecFN_small.scala 267:15]
  wire [2:0] divSqrtRecFNToRaw_io_roundingMode; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_io_rawOutValid_sqrt; // @[DivSqrtRecFN_small.scala 267:15]
  wire [2:0] divSqrtRecFNToRaw_io_roundingModeOut; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_io_invalidExc; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_io_infiniteExc; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_io_rawOut_sign; // @[DivSqrtRecFN_small.scala 267:15]
  wire [9:0] divSqrtRecFNToRaw_io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 267:15]
  wire [26:0] divSqrtRecFNToRaw_io_rawOut_sig; // @[DivSqrtRecFN_small.scala 267:15]
  wire [29:0] divSqrtRecFNToRaw_io_covSum; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_metaAssert; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_metaReset; // @[DivSqrtRecFN_small.scala 267:15]
  wire  roundRawFNToRecFN_io_invalidExc; // @[DivSqrtRecFN_small.scala 282:15]
  wire  roundRawFNToRecFN_io_infiniteExc; // @[DivSqrtRecFN_small.scala 282:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[DivSqrtRecFN_small.scala 282:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[DivSqrtRecFN_small.scala 282:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[DivSqrtRecFN_small.scala 282:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[DivSqrtRecFN_small.scala 282:15]
  wire [9:0] roundRawFNToRecFN_io_in_sExp; // @[DivSqrtRecFN_small.scala 282:15]
  wire [26:0] roundRawFNToRecFN_io_in_sig; // @[DivSqrtRecFN_small.scala 282:15]
  wire [2:0] roundRawFNToRecFN_io_roundingMode; // @[DivSqrtRecFN_small.scala 282:15]
  wire  roundRawFNToRecFN_io_detectTininess; // @[DivSqrtRecFN_small.scala 282:15]
  wire [32:0] roundRawFNToRecFN_io_out; // @[DivSqrtRecFN_small.scala 282:15]
  wire [4:0] roundRawFNToRecFN_io_exceptionFlags; // @[DivSqrtRecFN_small.scala 282:15]
  wire [29:0] roundRawFNToRecFN_io_covSum; // @[DivSqrtRecFN_small.scala 282:15]
  wire  roundRawFNToRecFN_metaAssert; // @[DivSqrtRecFN_small.scala 282:15]
  wire [29:0] DivSqrtRecFN_small_covSum;
  wire [29:0] divSqrtRecFNToRaw_sum;
  wire [29:0] roundRawFNToRecFN_sum;
  wire  divSqrtRecFNToRaw_metaAssert_wire;
  wire  roundRawFNToRecFN_metaAssert_wire;
  wire  DivSqrtRecFN_small_or0;
  reg  DivSqrtRecFN_small_metaAssert;
  reg [31:0] _RAND_0;
  DivSqrtRecFNToRaw_small divSqrtRecFNToRaw ( // @[DivSqrtRecFN_small.scala 267:15]
    .clock(divSqrtRecFNToRaw_clock),
    .reset(divSqrtRecFNToRaw_reset),
    .io_inReady(divSqrtRecFNToRaw_io_inReady),
    .io_inValid(divSqrtRecFNToRaw_io_inValid),
    .io_sqrtOp(divSqrtRecFNToRaw_io_sqrtOp),
    .io_a(divSqrtRecFNToRaw_io_a),
    .io_b(divSqrtRecFNToRaw_io_b),
    .io_roundingMode(divSqrtRecFNToRaw_io_roundingMode),
    .io_rawOutValid_div(divSqrtRecFNToRaw_io_rawOutValid_div),
    .io_rawOutValid_sqrt(divSqrtRecFNToRaw_io_rawOutValid_sqrt),
    .io_roundingModeOut(divSqrtRecFNToRaw_io_roundingModeOut),
    .io_invalidExc(divSqrtRecFNToRaw_io_invalidExc),
    .io_infiniteExc(divSqrtRecFNToRaw_io_infiniteExc),
    .io_rawOut_isNaN(divSqrtRecFNToRaw_io_rawOut_isNaN),
    .io_rawOut_isInf(divSqrtRecFNToRaw_io_rawOut_isInf),
    .io_rawOut_isZero(divSqrtRecFNToRaw_io_rawOut_isZero),
    .io_rawOut_sign(divSqrtRecFNToRaw_io_rawOut_sign),
    .io_rawOut_sExp(divSqrtRecFNToRaw_io_rawOut_sExp),
    .io_rawOut_sig(divSqrtRecFNToRaw_io_rawOut_sig),
    .io_covSum(divSqrtRecFNToRaw_io_covSum),
    .metaAssert(divSqrtRecFNToRaw_metaAssert),
    .metaReset(divSqrtRecFNToRaw_metaReset)
  );
  RoundRawFNToRecFN_2 roundRawFNToRecFN ( // @[DivSqrtRecFN_small.scala 282:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_infiniteExc(roundRawFNToRecFN_io_infiniteExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundRawFNToRecFN_io_detectTininess),
    .io_out(roundRawFNToRecFN_io_out),
    .io_exceptionFlags(roundRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundRawFNToRecFN_io_covSum),
    .metaAssert(roundRawFNToRecFN_metaAssert)
  );
  assign io_inReady = divSqrtRecFNToRaw_io_inReady; // @[DivSqrtRecFN_small.scala 269:16]
  assign io_outValid_div = divSqrtRecFNToRaw_io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 278:22]
  assign io_outValid_sqrt = divSqrtRecFNToRaw_io_rawOutValid_sqrt; // @[DivSqrtRecFN_small.scala 279:22]
  assign io_out = roundRawFNToRecFN_io_out; // @[DivSqrtRecFN_small.scala 288:23]
  assign io_exceptionFlags = roundRawFNToRecFN_io_exceptionFlags; // @[DivSqrtRecFN_small.scala 289:23]
  assign divSqrtRecFNToRaw_clock = clock;
  assign divSqrtRecFNToRaw_reset = reset;
  assign divSqrtRecFNToRaw_io_inValid = io_inValid; // @[DivSqrtRecFN_small.scala 270:39]
  assign divSqrtRecFNToRaw_io_sqrtOp = io_sqrtOp; // @[DivSqrtRecFN_small.scala 271:39]
  assign divSqrtRecFNToRaw_io_a = io_a; // @[DivSqrtRecFN_small.scala 272:39]
  assign divSqrtRecFNToRaw_io_b = io_b; // @[DivSqrtRecFN_small.scala 273:39]
  assign divSqrtRecFNToRaw_io_roundingMode = io_roundingMode; // @[DivSqrtRecFN_small.scala 274:39]
  assign roundRawFNToRecFN_io_invalidExc = divSqrtRecFNToRaw_io_invalidExc; // @[DivSqrtRecFN_small.scala 283:39]
  assign roundRawFNToRecFN_io_infiniteExc = divSqrtRecFNToRaw_io_infiniteExc; // @[DivSqrtRecFN_small.scala 284:39]
  assign roundRawFNToRecFN_io_in_isNaN = divSqrtRecFNToRaw_io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 285:39]
  assign roundRawFNToRecFN_io_in_isInf = divSqrtRecFNToRaw_io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 285:39]
  assign roundRawFNToRecFN_io_in_isZero = divSqrtRecFNToRaw_io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 285:39]
  assign roundRawFNToRecFN_io_in_sign = divSqrtRecFNToRaw_io_rawOut_sign; // @[DivSqrtRecFN_small.scala 285:39]
  assign roundRawFNToRecFN_io_in_sExp = divSqrtRecFNToRaw_io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 285:39]
  assign roundRawFNToRecFN_io_in_sig = divSqrtRecFNToRaw_io_rawOut_sig; // @[DivSqrtRecFN_small.scala 285:39]
  assign roundRawFNToRecFN_io_roundingMode = divSqrtRecFNToRaw_io_roundingModeOut; // @[DivSqrtRecFN_small.scala 286:39]
  assign roundRawFNToRecFN_io_detectTininess = 1'h1; // @[DivSqrtRecFN_small.scala 287:41]
  assign DivSqrtRecFN_small_covSum = 30'h0;
  assign divSqrtRecFNToRaw_sum = DivSqrtRecFN_small_covSum + divSqrtRecFNToRaw_io_covSum;
  assign roundRawFNToRecFN_sum = divSqrtRecFNToRaw_sum + roundRawFNToRecFN_io_covSum;
  assign io_covSum = roundRawFNToRecFN_sum;
  assign divSqrtRecFNToRaw_metaAssert_wire = divSqrtRecFNToRaw_metaAssert;
  assign roundRawFNToRecFN_metaAssert_wire = roundRawFNToRecFN_metaAssert;
  assign DivSqrtRecFN_small_or0 = divSqrtRecFNToRaw_metaAssert_wire | roundRawFNToRecFN_metaAssert_wire;
  assign metaAssert = DivSqrtRecFN_small_metaAssert;
  assign divSqrtRecFNToRaw_metaReset = metaReset | divSqrtRecFNToRaw_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  DivSqrtRecFN_small_metaAssert = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      DivSqrtRecFN_small_metaAssert <= 1'h0;
    end else begin
      DivSqrtRecFN_small_metaAssert <= DivSqrtRecFN_small_metaAssert | DivSqrtRecFN_small_or0;
    end
  end
endmodule
module DivSqrtRecFN_small_1(
  input         clock,
  input         reset,
  output        io_inReady,
  input         io_inValid,
  input         io_sqrtOp,
  input  [64:0] io_a,
  input  [64:0] io_b,
  input  [2:0]  io_roundingMode,
  output        io_outValid_div,
  output        io_outValid_sqrt,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         divSqrtRecFNToRaw_halt
);
  wire  divSqrtRecFNToRaw_clock; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_reset; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_io_inReady; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_io_inValid; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_io_sqrtOp; // @[DivSqrtRecFN_small.scala 267:15]
  wire [64:0] divSqrtRecFNToRaw_io_a; // @[DivSqrtRecFN_small.scala 267:15]
  wire [64:0] divSqrtRecFNToRaw_io_b; // @[DivSqrtRecFN_small.scala 267:15]
  wire [2:0] divSqrtRecFNToRaw_io_roundingMode; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_io_rawOutValid_sqrt; // @[DivSqrtRecFN_small.scala 267:15]
  wire [2:0] divSqrtRecFNToRaw_io_roundingModeOut; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_io_invalidExc; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_io_infiniteExc; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_io_rawOut_sign; // @[DivSqrtRecFN_small.scala 267:15]
  wire [12:0] divSqrtRecFNToRaw_io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 267:15]
  wire [55:0] divSqrtRecFNToRaw_io_rawOut_sig; // @[DivSqrtRecFN_small.scala 267:15]
  wire [29:0] divSqrtRecFNToRaw_io_covSum; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_metaAssert; // @[DivSqrtRecFN_small.scala 267:15]
  wire  divSqrtRecFNToRaw_metaReset; // @[DivSqrtRecFN_small.scala 267:15]
  wire  roundRawFNToRecFN_io_invalidExc; // @[DivSqrtRecFN_small.scala 282:15]
  wire  roundRawFNToRecFN_io_infiniteExc; // @[DivSqrtRecFN_small.scala 282:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[DivSqrtRecFN_small.scala 282:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[DivSqrtRecFN_small.scala 282:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[DivSqrtRecFN_small.scala 282:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[DivSqrtRecFN_small.scala 282:15]
  wire [12:0] roundRawFNToRecFN_io_in_sExp; // @[DivSqrtRecFN_small.scala 282:15]
  wire [55:0] roundRawFNToRecFN_io_in_sig; // @[DivSqrtRecFN_small.scala 282:15]
  wire [2:0] roundRawFNToRecFN_io_roundingMode; // @[DivSqrtRecFN_small.scala 282:15]
  wire  roundRawFNToRecFN_io_detectTininess; // @[DivSqrtRecFN_small.scala 282:15]
  wire [64:0] roundRawFNToRecFN_io_out; // @[DivSqrtRecFN_small.scala 282:15]
  wire [4:0] roundRawFNToRecFN_io_exceptionFlags; // @[DivSqrtRecFN_small.scala 282:15]
  wire [29:0] roundRawFNToRecFN_io_covSum; // @[DivSqrtRecFN_small.scala 282:15]
  wire  roundRawFNToRecFN_metaAssert; // @[DivSqrtRecFN_small.scala 282:15]
  wire [29:0] DivSqrtRecFN_small_1_covSum;
  wire [29:0] divSqrtRecFNToRaw_sum;
  wire [29:0] roundRawFNToRecFN_sum;
  wire  divSqrtRecFNToRaw_metaAssert_wire;
  wire  roundRawFNToRecFN_metaAssert_wire;
  wire  DivSqrtRecFN_small_1_or0;
  reg  DivSqrtRecFN_small_1_metaAssert;
  reg [31:0] _RAND_0;
  DivSqrtRecFNToRaw_small_1 divSqrtRecFNToRaw ( // @[DivSqrtRecFN_small.scala 267:15]
    .clock(divSqrtRecFNToRaw_clock),
    .reset(divSqrtRecFNToRaw_reset),
    .io_inReady(divSqrtRecFNToRaw_io_inReady),
    .io_inValid(divSqrtRecFNToRaw_io_inValid),
    .io_sqrtOp(divSqrtRecFNToRaw_io_sqrtOp),
    .io_a(divSqrtRecFNToRaw_io_a),
    .io_b(divSqrtRecFNToRaw_io_b),
    .io_roundingMode(divSqrtRecFNToRaw_io_roundingMode),
    .io_rawOutValid_div(divSqrtRecFNToRaw_io_rawOutValid_div),
    .io_rawOutValid_sqrt(divSqrtRecFNToRaw_io_rawOutValid_sqrt),
    .io_roundingModeOut(divSqrtRecFNToRaw_io_roundingModeOut),
    .io_invalidExc(divSqrtRecFNToRaw_io_invalidExc),
    .io_infiniteExc(divSqrtRecFNToRaw_io_infiniteExc),
    .io_rawOut_isNaN(divSqrtRecFNToRaw_io_rawOut_isNaN),
    .io_rawOut_isInf(divSqrtRecFNToRaw_io_rawOut_isInf),
    .io_rawOut_isZero(divSqrtRecFNToRaw_io_rawOut_isZero),
    .io_rawOut_sign(divSqrtRecFNToRaw_io_rawOut_sign),
    .io_rawOut_sExp(divSqrtRecFNToRaw_io_rawOut_sExp),
    .io_rawOut_sig(divSqrtRecFNToRaw_io_rawOut_sig),
    .io_covSum(divSqrtRecFNToRaw_io_covSum),
    .metaAssert(divSqrtRecFNToRaw_metaAssert),
    .metaReset(divSqrtRecFNToRaw_metaReset)
  );
  RoundRawFNToRecFN_3 roundRawFNToRecFN ( // @[DivSqrtRecFN_small.scala 282:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_infiniteExc(roundRawFNToRecFN_io_infiniteExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundRawFNToRecFN_io_detectTininess),
    .io_out(roundRawFNToRecFN_io_out),
    .io_exceptionFlags(roundRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundRawFNToRecFN_io_covSum),
    .metaAssert(roundRawFNToRecFN_metaAssert)
  );
  assign io_inReady = divSqrtRecFNToRaw_io_inReady; // @[DivSqrtRecFN_small.scala 269:16]
  assign io_outValid_div = divSqrtRecFNToRaw_io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 278:22]
  assign io_outValid_sqrt = divSqrtRecFNToRaw_io_rawOutValid_sqrt; // @[DivSqrtRecFN_small.scala 279:22]
  assign io_out = roundRawFNToRecFN_io_out; // @[DivSqrtRecFN_small.scala 288:23]
  assign io_exceptionFlags = roundRawFNToRecFN_io_exceptionFlags; // @[DivSqrtRecFN_small.scala 289:23]
  assign divSqrtRecFNToRaw_clock = clock;
  assign divSqrtRecFNToRaw_reset = reset;
  assign divSqrtRecFNToRaw_io_inValid = io_inValid; // @[DivSqrtRecFN_small.scala 270:39]
  assign divSqrtRecFNToRaw_io_sqrtOp = io_sqrtOp; // @[DivSqrtRecFN_small.scala 271:39]
  assign divSqrtRecFNToRaw_io_a = io_a; // @[DivSqrtRecFN_small.scala 272:39]
  assign divSqrtRecFNToRaw_io_b = io_b; // @[DivSqrtRecFN_small.scala 273:39]
  assign divSqrtRecFNToRaw_io_roundingMode = io_roundingMode; // @[DivSqrtRecFN_small.scala 274:39]
  assign roundRawFNToRecFN_io_invalidExc = divSqrtRecFNToRaw_io_invalidExc; // @[DivSqrtRecFN_small.scala 283:39]
  assign roundRawFNToRecFN_io_infiniteExc = divSqrtRecFNToRaw_io_infiniteExc; // @[DivSqrtRecFN_small.scala 284:39]
  assign roundRawFNToRecFN_io_in_isNaN = divSqrtRecFNToRaw_io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 285:39]
  assign roundRawFNToRecFN_io_in_isInf = divSqrtRecFNToRaw_io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 285:39]
  assign roundRawFNToRecFN_io_in_isZero = divSqrtRecFNToRaw_io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 285:39]
  assign roundRawFNToRecFN_io_in_sign = divSqrtRecFNToRaw_io_rawOut_sign; // @[DivSqrtRecFN_small.scala 285:39]
  assign roundRawFNToRecFN_io_in_sExp = divSqrtRecFNToRaw_io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 285:39]
  assign roundRawFNToRecFN_io_in_sig = divSqrtRecFNToRaw_io_rawOut_sig; // @[DivSqrtRecFN_small.scala 285:39]
  assign roundRawFNToRecFN_io_roundingMode = divSqrtRecFNToRaw_io_roundingModeOut; // @[DivSqrtRecFN_small.scala 286:39]
  assign roundRawFNToRecFN_io_detectTininess = 1'h1; // @[DivSqrtRecFN_small.scala 287:41]
  assign DivSqrtRecFN_small_1_covSum = 30'h0;
  assign divSqrtRecFNToRaw_sum = DivSqrtRecFN_small_1_covSum + divSqrtRecFNToRaw_io_covSum;
  assign roundRawFNToRecFN_sum = divSqrtRecFNToRaw_sum + roundRawFNToRecFN_io_covSum;
  assign io_covSum = roundRawFNToRecFN_sum;
  assign divSqrtRecFNToRaw_metaAssert_wire = divSqrtRecFNToRaw_metaAssert;
  assign roundRawFNToRecFN_metaAssert_wire = roundRawFNToRecFN_metaAssert;
  assign DivSqrtRecFN_small_1_or0 = divSqrtRecFNToRaw_metaAssert_wire | roundRawFNToRecFN_metaAssert_wire;
  assign metaAssert = DivSqrtRecFN_small_1_metaAssert;
  assign divSqrtRecFNToRaw_metaReset = metaReset | divSqrtRecFNToRaw_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  DivSqrtRecFN_small_1_metaAssert = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      DivSqrtRecFN_small_1_metaAssert <= 1'h0;
    end else begin
      DivSqrtRecFN_small_1_metaAssert <= DivSqrtRecFN_small_1_metaAssert | DivSqrtRecFN_small_1_or0;
    end
  end
endmodule
module RRArbiter(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [26:0] io_in_0_bits_bits_addr,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input         io_in_1_bits_valid,
  input  [26:0] io_in_1_bits_bits_addr,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_valid,
  output [26:0] io_out_bits_bits_addr,
  output        io_chosen,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire  _T_104; // @[Decoupled.scala 37:37]
  reg  _T_106; // @[Reg.scala 11:16]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[Arbiter.scala 67:57]
  wire  _T_110; // @[Arbiter.scala 68:83]
  wire  _T_112; // @[Arbiter.scala 31:68]
  wire  _T_119; // @[Arbiter.scala 72:50]
  wire  _GEN_9; // @[Arbiter.scala 77:27]
  wire [29:0] RRArbiter_covSum;
  assign _T_104 = io_out_ready & io_out_valid; // @[Decoupled.scala 37:37]
  assign _T_108 = 1'h1 > _T_106; // @[Arbiter.scala 67:57]
  assign _T_110 = io_in_1_valid & _T_108; // @[Arbiter.scala 68:83]
  assign _T_112 = _T_110 | io_in_0_valid; // @[Arbiter.scala 31:68]
  assign _T_119 = _T_108 | ~_T_112; // @[Arbiter.scala 72:50]
  assign _GEN_9 = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 77:27]
  assign io_in_0_ready = ~_T_110 & io_out_ready; // @[Arbiter.scala 60:16]
  assign io_in_1_ready = _T_119 & io_out_ready; // @[Arbiter.scala 60:16]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16]
  assign io_out_bits_valid = io_chosen ? io_in_1_bits_valid : 1'h1; // @[Arbiter.scala 42:15]
  assign io_out_bits_bits_addr = io_chosen ? io_in_1_bits_bits_addr : io_in_0_bits_bits_addr; // @[Arbiter.scala 42:15]
  assign io_chosen = _T_110 | _GEN_9; // @[Arbiter.scala 40:13]
  assign RRArbiter_covSum = 30'h0;
  assign io_covSum = RRArbiter_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_106 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      _T_106 <= 1'h0;
    end else if (_T_104) begin
      _T_106 <= io_chosen;
    end
  end
endmodule
module PCodeLock(
  input  [53:0] io_in_ppn,
  input  [1:0]  io_in_reserved_for_software,
  input         io_in_d,
  input         io_in_a,
  input         io_in_g,
  input         io_in_u,
  input         io_in_x,
  input         io_in_w,
  input         io_in_r,
  input         io_in_v,
  output [53:0] io_out_ppn,
  output [1:0]  io_out_reserved_for_software,
  output        io_out_d,
  output        io_out_a,
  output        io_out_g,
  output        io_out_u,
  output        io_out_x,
  output        io_out_w,
  output        io_out_r,
  output        io_out_v,
  input  [19:0] io_cfg_0_base,
  input  [9:0]  io_cfg_0_mask,
  input         io_cfg_0_valid,
  input         io_cfg_0_enable,
  input  [19:0] io_cfg_1_base,
  input  [9:0]  io_cfg_1_mask,
  input         io_cfg_1_valid,
  input         io_cfg_1_enable,
  input  [19:0] io_cfg_2_base,
  input  [9:0]  io_cfg_2_mask,
  input         io_cfg_2_valid,
  input         io_cfg_2_enable,
  input  [19:0] io_cfg_3_base,
  input  [9:0]  io_cfg_3_mask,
  input         io_cfg_3_valid,
  input         io_cfg_3_enable,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  _T_16; // @[PTW.scala 108:58]
  wire  _T_17; // @[PTW.scala 108:58]
  wire  enable; // @[PTW.scala 108:58]
  wire  _T_20; // @[PTW.scala 77:44]
  wire  _T_21; // @[PTW.scala 77:38]
  wire  _T_22; // @[PTW.scala 77:32]
  wire  _T_23; // @[PTW.scala 77:52]
  wire  _T_25; // @[PTW.scala 124:26]
  wire  _T_26; // @[PTW.scala 127:28]
  wire [19:0] _T_28; // @[Cat.scala 30:58]
  wire [19:0] _T_30; // @[PTW.scala 114:72]
  wire  _T_31; // @[PTW.scala 114:101]
  wire  _T_32; // @[PTW.scala 114:20]
  wire [19:0] _T_34; // @[Cat.scala 30:58]
  wire [19:0] _T_36; // @[PTW.scala 114:72]
  wire  _T_37; // @[PTW.scala 114:101]
  wire  _T_38; // @[PTW.scala 114:20]
  wire [19:0] _T_40; // @[Cat.scala 30:58]
  wire [19:0] _T_42; // @[PTW.scala 114:72]
  wire  _T_43; // @[PTW.scala 114:101]
  wire  _T_44; // @[PTW.scala 114:20]
  wire [19:0] _T_46; // @[Cat.scala 30:58]
  wire [19:0] _T_48; // @[PTW.scala 114:72]
  wire  _T_49; // @[PTW.scala 114:101]
  wire  _T_50; // @[PTW.scala 114:20]
  wire  _T_52; // @[PTW.scala 115:49]
  wire  _T_53; // @[PTW.scala 115:49]
  wire  _T_54; // @[PTW.scala 115:49]
  wire  _T_93; // @[PTW.scala 128:41]
  wire [29:0] PCodeLock_covSum;
  assign _T_16 = io_cfg_0_enable & io_cfg_1_enable; // @[PTW.scala 108:58]
  assign _T_17 = _T_16 & io_cfg_2_enable; // @[PTW.scala 108:58]
  assign enable = _T_17 & io_cfg_3_enable; // @[PTW.scala 108:58]
  assign _T_20 = io_in_x & ~io_in_w; // @[PTW.scala 77:44]
  assign _T_21 = io_in_r | _T_20; // @[PTW.scala 77:38]
  assign _T_22 = io_in_v & _T_21; // @[PTW.scala 77:32]
  assign _T_23 = _T_22 & io_in_a; // @[PTW.scala 77:52]
  assign _T_25 = ~enable | ~_T_23; // @[PTW.scala 124:26]
  assign _T_26 = _T_25 | io_in_u; // @[PTW.scala 127:28]
  assign _T_28 = {8'hff,io_cfg_0_mask,2'h0}; // @[Cat.scala 30:58]
  assign _T_30 = _T_28 & io_in_ppn[19:0]; // @[PTW.scala 114:72]
  assign _T_31 = _T_30 == io_cfg_0_base; // @[PTW.scala 114:101]
  assign _T_32 = io_cfg_0_valid & _T_31; // @[PTW.scala 114:20]
  assign _T_34 = {8'hff,io_cfg_1_mask,2'h0}; // @[Cat.scala 30:58]
  assign _T_36 = _T_34 & io_in_ppn[19:0]; // @[PTW.scala 114:72]
  assign _T_37 = _T_36 == io_cfg_1_base; // @[PTW.scala 114:101]
  assign _T_38 = io_cfg_1_valid & _T_37; // @[PTW.scala 114:20]
  assign _T_40 = {8'hff,io_cfg_2_mask,2'h0}; // @[Cat.scala 30:58]
  assign _T_42 = _T_40 & io_in_ppn[19:0]; // @[PTW.scala 114:72]
  assign _T_43 = _T_42 == io_cfg_2_base; // @[PTW.scala 114:101]
  assign _T_44 = io_cfg_2_valid & _T_43; // @[PTW.scala 114:20]
  assign _T_46 = {8'hff,io_cfg_3_mask,2'h0}; // @[Cat.scala 30:58]
  assign _T_48 = _T_46 & io_in_ppn[19:0]; // @[PTW.scala 114:72]
  assign _T_49 = _T_48 == io_cfg_3_base; // @[PTW.scala 114:101]
  assign _T_50 = io_cfg_3_valid & _T_49; // @[PTW.scala 114:20]
  assign _T_52 = _T_32 | _T_38; // @[PTW.scala 115:49]
  assign _T_53 = _T_52 | _T_44; // @[PTW.scala 115:49]
  assign _T_54 = _T_53 | _T_50; // @[PTW.scala 115:49]
  assign _T_93 = _T_54 ? 1'h0 : io_in_w; // @[PTW.scala 128:41]
  assign io_out_ppn = io_in_ppn; // @[PTW.scala 106:12]
  assign io_out_reserved_for_software = io_in_reserved_for_software; // @[PTW.scala 106:12]
  assign io_out_d = io_in_d; // @[PTW.scala 106:12]
  assign io_out_a = io_in_a; // @[PTW.scala 106:12]
  assign io_out_g = io_in_g; // @[PTW.scala 106:12]
  assign io_out_u = io_in_u; // @[PTW.scala 106:12]
  assign io_out_x = _T_26 ? io_in_x : _T_54; // @[PTW.scala 106:12 PTW.scala 127:14]
  assign io_out_w = _T_25 ? io_in_w : _T_93; // @[PTW.scala 106:12 PTW.scala 128:14]
  assign io_out_r = io_in_r; // @[PTW.scala 106:12]
  assign io_out_v = io_in_v; // @[PTW.scala 106:12]
  assign PCodeLock_covSum = 30'h0;
  assign io_covSum = PCodeLock_covSum;
  assign metaAssert = 1'h0;
endmodule
module IBuf(
  input         clock,
  input         reset,
  output        io_imem_ready,
  input         io_imem_valid,
  input         io_imem_bits_btb_taken,
  input         io_imem_bits_btb_bridx,
  input  [4:0]  io_imem_bits_btb_entry,
  input  [7:0]  io_imem_bits_btb_bht_history,
  input  [39:0] io_imem_bits_pc,
  input  [31:0] io_imem_bits_data,
  input         io_imem_bits_xcpt_pf_inst,
  input         io_imem_bits_xcpt_ae_inst,
  input         io_imem_bits_replay,
  input         io_kill,
  output [39:0] io_pc,
  output [4:0]  io_btb_resp_entry,
  output [7:0]  io_btb_resp_bht_history,
  input         io_inst_0_ready,
  output        io_inst_0_valid,
  output        io_inst_0_bits_xcpt0_pf_inst,
  output        io_inst_0_bits_xcpt0_ae_inst,
  output        io_inst_0_bits_xcpt1_pf_inst,
  output        io_inst_0_bits_xcpt1_ae_inst,
  output        io_inst_0_bits_replay,
  output        io_inst_0_bits_rvc,
  output [31:0] io_inst_0_bits_inst_bits,
  output [4:0]  io_inst_0_bits_inst_rd,
  output [4:0]  io_inst_0_bits_inst_rs1,
  output [4:0]  io_inst_0_bits_inst_rs2,
  output [4:0]  io_inst_0_bits_inst_rs3,
  output [31:0] io_inst_0_bits_raw,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [31:0] RVCExpander_io_in; // @[IBuf.scala 86:21]
  wire [31:0] RVCExpander_io_out_bits; // @[IBuf.scala 86:21]
  wire [4:0] RVCExpander_io_out_rd; // @[IBuf.scala 86:21]
  wire [4:0] RVCExpander_io_out_rs1; // @[IBuf.scala 86:21]
  wire [4:0] RVCExpander_io_out_rs2; // @[IBuf.scala 86:21]
  wire [4:0] RVCExpander_io_out_rs3; // @[IBuf.scala 86:21]
  wire  RVCExpander_io_rvc; // @[IBuf.scala 86:21]
  wire [29:0] RVCExpander_io_covSum; // @[IBuf.scala 86:21]
  wire  RVCExpander_metaAssert; // @[IBuf.scala 86:21]
  reg  nBufValid; // @[IBuf.scala 34:47]
  reg [31:0] _RAND_0;
  reg [39:0] buf__pc; // @[IBuf.scala 35:16]
  reg [63:0] _RAND_1;
  reg [31:0] buf__data; // @[IBuf.scala 35:16]
  reg [31:0] _RAND_2;
  reg  buf__xcpt_pf_inst; // @[IBuf.scala 35:16]
  reg [31:0] _RAND_3;
  reg  buf__xcpt_ae_inst; // @[IBuf.scala 35:16]
  reg [31:0] _RAND_4;
  reg  buf__replay; // @[IBuf.scala 35:16]
  reg [31:0] _RAND_5;
  reg [4:0] ibufBTBResp_entry; // @[IBuf.scala 36:24]
  reg [31:0] _RAND_6;
  reg [7:0] ibufBTBResp_bht_history; // @[IBuf.scala 36:24]
  reg [31:0] _RAND_7;
  wire  pcWordBits; // @[package.scala 119:13]
  wire [1:0] _T_25; // @[IBuf.scala 41:64]
  wire [1:0] _T_26; // @[IBuf.scala 41:16]
  wire [1:0] _GEN_56; // @[IBuf.scala 41:88]
  wire [1:0] nIC; // @[IBuf.scala 41:88]
  wire [1:0] _T_31; // @[IBuf.scala 43:19]
  wire [1:0] _GEN_57; // @[IBuf.scala 43:49]
  wire [1:0] nValid; // @[IBuf.scala 43:49]
  wire [3:0] _T_94; // @[OneHot.scala 45:35]
  wire [3:0] _T_97; // @[IBuf.scala 74:33]
  wire [1:0] valid; // @[IBuf.scala 74:37]
  wire [1:0] _T_127; // @[IBuf.scala 93:42]
  wire  _T_129; // @[IBuf.scala 93:34]
  wire [1:0] _T_98; // @[OneHot.scala 45:35]
  wire [1:0] bufMask; // @[IBuf.scala 75:37]
  wire [1:0] buf_replay; // @[IBuf.scala 77:23]
  wire  _T_132; // @[IBuf.scala 93:48]
  wire [1:0] _T_165; // @[IBuf.scala 102:71]
  wire [1:0] nReady; // @[IBuf.scala 102:56]
  wire [1:0] nICReady; // @[IBuf.scala 42:25]
  wire  _T_33; // @[IBuf.scala 44:47]
  wire  _T_34; // @[IBuf.scala 44:37]
  wire  _T_35; // @[IBuf.scala 44:73]
  wire [1:0] _T_38; // @[IBuf.scala 44:92]
  wire  _T_39; // @[IBuf.scala 44:85]
  wire  _T_40; // @[IBuf.scala 44:80]
  wire [1:0] _T_45; // @[IBuf.scala 48:64]
  wire [1:0] _T_46; // @[IBuf.scala 48:23]
  wire  _T_48; // @[IBuf.scala 54:27]
  wire  _T_49; // @[IBuf.scala 54:62]
  wire  _T_50; // @[IBuf.scala 54:50]
  wire  _T_55; // @[IBuf.scala 54:68]
  wire [1:0] _T_57; // @[IBuf.scala 55:32]
  wire [63:0] _T_63; // @[Cat.scala 30:58]
  wire [5:0] _T_64; // @[IBuf.scala 128:19]
  wire [63:0] _T_65; // @[IBuf.scala 128:10]
  wire [39:0] _T_68; // @[IBuf.scala 59:35]
  wire [2:0] _T_69; // @[IBuf.scala 59:80]
  wire [39:0] _GEN_65; // @[IBuf.scala 59:68]
  wire [39:0] _T_71; // @[IBuf.scala 59:68]
  wire [39:0] _T_72; // @[IBuf.scala 59:109]
  wire [39:0] _T_73; // @[IBuf.scala 59:49]
  wire [1:0] _GEN_0; // @[IBuf.scala 54:92]
  wire [1:0] _GEN_23; // @[IBuf.scala 47:29]
  wire [1:0] _GEN_46; // @[IBuf.scala 63:20]
  wire [1:0] _T_75; // @[IBuf.scala 68:32]
  wire [1:0] icShiftAmt; // @[IBuf.scala 68:44]
  wire [63:0] _T_81; // @[Cat.scala 30:58]
  wire [127:0] _T_85; // @[Cat.scala 30:58]
  wire [5:0] _T_86; // @[IBuf.scala 121:19]
  wire [190:0] _GEN_68; // @[IBuf.scala 121:10]
  wire [190:0] _T_87; // @[IBuf.scala 121:10]
  wire [31:0] icData; // @[package.scala 119:13]
  wire [4:0] _T_89; // @[IBuf.scala 71:65]
  wire [62:0] _T_90; // @[IBuf.scala 71:51]
  wire [31:0] icMask; // @[IBuf.scala 71:92]
  wire [31:0] _T_91; // @[IBuf.scala 72:21]
  wire [31:0] _T_93; // @[IBuf.scala 72:41]
  wire  xcpt_1_pf_inst; // @[IBuf.scala 76:53]
  wire  xcpt_1_ae_inst; // @[IBuf.scala 76:53]
  wire [1:0] _T_104; // @[IBuf.scala 78:63]
  wire [1:0] _T_105; // @[IBuf.scala 78:35]
  wire [1:0] ic_replay; // @[IBuf.scala 78:30]
  wire  _T_108; // @[IBuf.scala 79:25]
  wire  _T_109; // @[IBuf.scala 79:78]
  wire  _T_110; // @[IBuf.scala 79:52]
  wire  _T_112; // @[IBuf.scala 79:9]
  wire  _T_114; // @[IBuf.scala 82:26]
  wire [1:0] _T_121; // @[IBuf.scala 92:61]
  wire  _T_123; // @[IBuf.scala 92:49]
  wire [1:0] _T_142; // @[IBuf.scala 96:63]
  wire [1:0] _T_143; // @[IBuf.scala 96:35]
  wire  _T_153; // @[IBuf.scala 100:25]
  wire [1:0] _T_156; // @[IBuf.scala 100:50]
  wire  _T_158; // @[IBuf.scala 100:40]
  reg [1:0] IBuf_state; // @[Register tracking IBuf state]
  reg [31:0] _RAND_8;
  reg  IBuf_cov [0:3]; // @[Coverage map for IBuf]
  reg [31:0] _RAND_9;
  wire  IBuf_cov_read_data; // @[Coverage map for IBuf]
  wire [1:0] IBuf_cov_read_addr; // @[Coverage map for IBuf]
  wire  IBuf_cov_write_data; // @[Coverage map for IBuf]
  wire [1:0] IBuf_cov_write_addr; // @[Coverage map for IBuf]
  wire  IBuf_cov_write_mask; // @[Coverage map for IBuf]
  wire  IBuf_cov_write_en; // @[Coverage map for IBuf]
  reg [29:0] IBuf_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_10;
  wire  nBufValid_shl;
  wire [1:0] nBufValid_pad;
  wire [1:0] buf__replay_shl;
  wire [1:0] buf__replay_pad;
  wire [1:0] IBuf_xor0;
  wire [29:0] RVCExpander_sum;
  wire  stopEn0;
  wire  RVCExpander_metaAssert_wire;
  wire  IBuf_or0;
  reg  IBuf_metaAssert;
  reg [31:0] _RAND_11;
  RVCExpander RVCExpander ( // @[IBuf.scala 86:21]
    .io_in(RVCExpander_io_in),
    .io_out_bits(RVCExpander_io_out_bits),
    .io_out_rd(RVCExpander_io_out_rd),
    .io_out_rs1(RVCExpander_io_out_rs1),
    .io_out_rs2(RVCExpander_io_out_rs2),
    .io_out_rs3(RVCExpander_io_out_rs3),
    .io_rvc(RVCExpander_io_rvc),
    .io_covSum(RVCExpander_io_covSum),
    .metaAssert(RVCExpander_metaAssert)
  );
  assign pcWordBits = io_imem_bits_pc[1]; // @[package.scala 119:13]
  assign _T_25 = io_imem_bits_btb_bridx + 1'h1; // @[IBuf.scala 41:64]
  assign _T_26 = io_imem_bits_btb_taken ? _T_25 : 2'h2; // @[IBuf.scala 41:16]
  assign _GEN_56 = {{1'd0}, pcWordBits}; // @[IBuf.scala 41:88]
  assign nIC = _T_26 - _GEN_56; // @[IBuf.scala 41:88]
  assign _T_31 = io_imem_valid ? nIC : 2'h0; // @[IBuf.scala 43:19]
  assign _GEN_57 = {{1'd0}, nBufValid}; // @[IBuf.scala 43:49]
  assign nValid = _T_31 + _GEN_57; // @[IBuf.scala 43:49]
  assign _T_94 = 4'h1 << nValid; // @[OneHot.scala 45:35]
  assign _T_97 = _T_94 - 4'h1; // @[IBuf.scala 74:33]
  assign valid = _T_97[1:0]; // @[IBuf.scala 74:37]
  assign _T_127 = {{1'd0}, valid[1]}; // @[IBuf.scala 93:42]
  assign _T_129 = RVCExpander_io_rvc | _T_127[0]; // @[IBuf.scala 93:34]
  assign _T_98 = 2'h1 << nBufValid; // @[OneHot.scala 45:35]
  assign bufMask = _T_98 - 2'h1; // @[IBuf.scala 75:37]
  assign buf_replay = buf__replay ? bufMask : 2'h0; // @[IBuf.scala 77:23]
  assign _T_132 = _T_129 | buf_replay[0]; // @[IBuf.scala 93:48]
  assign _T_165 = RVCExpander_io_rvc ? 2'h1 : 2'h2; // @[IBuf.scala 102:71]
  assign nReady = _T_132 ? _T_165 : 2'h0; // @[IBuf.scala 102:56]
  assign nICReady = nReady - _GEN_57; // @[IBuf.scala 42:25]
  assign _T_33 = nReady >= _GEN_57; // @[IBuf.scala 44:47]
  assign _T_34 = io_inst_0_ready & _T_33; // @[IBuf.scala 44:37]
  assign _T_35 = nICReady >= nIC; // @[IBuf.scala 44:73]
  assign _T_38 = nIC - nICReady; // @[IBuf.scala 44:92]
  assign _T_39 = 2'h1 >= _T_38; // @[IBuf.scala 44:85]
  assign _T_40 = _T_35 | _T_39; // @[IBuf.scala 44:80]
  assign _T_45 = _GEN_57 - nReady; // @[IBuf.scala 48:64]
  assign _T_46 = _T_33 ? 2'h0 : _T_45; // @[IBuf.scala 48:23]
  assign _T_48 = io_imem_valid & _T_33; // @[IBuf.scala 54:27]
  assign _T_49 = nICReady < nIC; // @[IBuf.scala 54:62]
  assign _T_50 = _T_48 & _T_49; // @[IBuf.scala 54:50]
  assign _T_55 = _T_50 & _T_39; // @[IBuf.scala 54:68]
  assign _T_57 = _GEN_56 + nICReady; // @[IBuf.scala 55:32]
  assign _T_63 = {io_imem_bits_data[31:16],io_imem_bits_data[31:16],io_imem_bits_data}; // @[Cat.scala 30:58]
  assign _T_64 = {_T_57, 4'h0}; // @[IBuf.scala 128:19]
  assign _T_65 = _T_63 >> _T_64; // @[IBuf.scala 128:10]
  assign _T_68 = io_imem_bits_pc & 40'hfffffffffc; // @[IBuf.scala 59:35]
  assign _T_69 = {nICReady, 1'h0}; // @[IBuf.scala 59:80]
  assign _GEN_65 = {{37'd0}, _T_69}; // @[IBuf.scala 59:68]
  assign _T_71 = io_imem_bits_pc + _GEN_65; // @[IBuf.scala 59:68]
  assign _T_72 = _T_71 & 40'h3; // @[IBuf.scala 59:109]
  assign _T_73 = _T_68 | _T_72; // @[IBuf.scala 59:49]
  assign _GEN_0 = _T_55 ? _T_38 : _T_46; // @[IBuf.scala 54:92]
  assign _GEN_23 = io_inst_0_ready ? _GEN_0 : {{1'd0}, nBufValid}; // @[IBuf.scala 47:29]
  assign _GEN_46 = io_kill ? 2'h0 : _GEN_23; // @[IBuf.scala 63:20]
  assign _T_75 = 2'h2 + _GEN_57; // @[IBuf.scala 68:32]
  assign icShiftAmt = _T_75 - _GEN_56; // @[IBuf.scala 68:44]
  assign _T_81 = {io_imem_bits_data,io_imem_bits_data[15:0],io_imem_bits_data[15:0]}; // @[Cat.scala 30:58]
  assign _T_85 = {_T_81[63:48],_T_81[63:48],_T_81[63:48],_T_81[63:48],io_imem_bits_data,io_imem_bits_data[15:0],io_imem_bits_data[15:0]}; // @[Cat.scala 30:58]
  assign _T_86 = {icShiftAmt, 4'h0}; // @[IBuf.scala 121:19]
  assign _GEN_68 = {{63'd0}, _T_85}; // @[IBuf.scala 121:10]
  assign _T_87 = _GEN_68 << _T_86; // @[IBuf.scala 121:10]
  assign icData = _T_87[95:64]; // @[package.scala 119:13]
  assign _T_89 = {nBufValid, 4'h0}; // @[IBuf.scala 71:65]
  assign _T_90 = 63'hffffffff << _T_89; // @[IBuf.scala 71:51]
  assign icMask = _T_90[31:0]; // @[IBuf.scala 71:92]
  assign _T_91 = icData & icMask; // @[IBuf.scala 72:21]
  assign _T_93 = buf__data & ~icMask; // @[IBuf.scala 72:41]
  assign xcpt_1_pf_inst = bufMask[1] ? buf__xcpt_pf_inst : io_imem_bits_xcpt_pf_inst; // @[IBuf.scala 76:53]
  assign xcpt_1_ae_inst = bufMask[1] ? buf__xcpt_ae_inst : io_imem_bits_xcpt_ae_inst; // @[IBuf.scala 76:53]
  assign _T_104 = valid & ~bufMask; // @[IBuf.scala 78:63]
  assign _T_105 = io_imem_bits_replay ? _T_104 : 2'h0; // @[IBuf.scala 78:35]
  assign ic_replay = buf_replay | _T_105; // @[IBuf.scala 78:30]
  assign _T_108 = ~io_imem_valid | ~io_imem_bits_btb_taken; // @[IBuf.scala 79:25]
  assign _T_109 = io_imem_bits_btb_bridx >= pcWordBits; // @[IBuf.scala 79:78]
  assign _T_110 = _T_108 | _T_109; // @[IBuf.scala 79:52]
  assign _T_112 = _T_110 | reset; // @[IBuf.scala 79:9]
  assign _T_114 = nBufValid > 1'h0; // @[IBuf.scala 82:26]
  assign _T_121 = {{1'd0}, ic_replay[1]}; // @[IBuf.scala 92:61]
  assign _T_123 = ~RVCExpander_io_rvc & _T_121[0]; // @[IBuf.scala 92:49]
  assign _T_142 = {xcpt_1_pf_inst,xcpt_1_ae_inst}; // @[IBuf.scala 96:63]
  assign _T_143 = RVCExpander_io_rvc ? 2'h0 : _T_142; // @[IBuf.scala 96:35]
  assign _T_153 = bufMask[0] & RVCExpander_io_rvc; // @[IBuf.scala 100:25]
  assign _T_156 = {{1'd0}, bufMask[1]}; // @[IBuf.scala 100:50]
  assign _T_158 = _T_153 | _T_156[0]; // @[IBuf.scala 100:40]
  assign io_imem_ready = _T_34 & _T_40; // @[IBuf.scala 44:17]
  assign io_pc = _T_114 ? buf__pc : io_imem_bits_pc; // @[IBuf.scala 82:9]
  assign io_btb_resp_entry = _T_158 ? ibufBTBResp_entry : io_imem_bits_btb_entry; // @[IBuf.scala 81:15 IBuf.scala 100:71]
  assign io_btb_resp_bht_history = _T_158 ? ibufBTBResp_bht_history : io_imem_bits_btb_bht_history; // @[IBuf.scala 81:15 IBuf.scala 100:71]
  assign io_inst_0_valid = valid[0] & _T_132; // @[IBuf.scala 94:24]
  assign io_inst_0_bits_xcpt0_pf_inst = bufMask[0] ? buf__xcpt_pf_inst : io_imem_bits_xcpt_pf_inst; // @[IBuf.scala 95:29]
  assign io_inst_0_bits_xcpt0_ae_inst = bufMask[0] ? buf__xcpt_ae_inst : io_imem_bits_xcpt_ae_inst; // @[IBuf.scala 95:29]
  assign io_inst_0_bits_xcpt1_pf_inst = _T_143[1]; // @[IBuf.scala 96:29]
  assign io_inst_0_bits_xcpt1_ae_inst = _T_143[0]; // @[IBuf.scala 96:29]
  assign io_inst_0_bits_replay = ic_replay[0] | _T_123; // @[IBuf.scala 97:30]
  assign io_inst_0_bits_rvc = RVCExpander_io_rvc; // @[IBuf.scala 98:27]
  assign io_inst_0_bits_inst_bits = RVCExpander_io_out_bits; // @[IBuf.scala 88:26]
  assign io_inst_0_bits_inst_rd = RVCExpander_io_out_rd; // @[IBuf.scala 88:26]
  assign io_inst_0_bits_inst_rs1 = RVCExpander_io_out_rs1; // @[IBuf.scala 88:26]
  assign io_inst_0_bits_inst_rs2 = RVCExpander_io_out_rs2; // @[IBuf.scala 88:26]
  assign io_inst_0_bits_inst_rs3 = RVCExpander_io_out_rs3; // @[IBuf.scala 88:26]
  assign io_inst_0_bits_raw = _T_91 | _T_93; // @[IBuf.scala 89:25]
  assign RVCExpander_io_in = _T_91 | _T_93; // @[IBuf.scala 87:15]
  assign IBuf_cov_read_addr = IBuf_state;
  assign IBuf_cov_read_data = IBuf_cov[IBuf_cov_read_addr]; // @[Coverage map for IBuf]
  assign IBuf_cov_write_data = 1'h1;
  assign IBuf_cov_write_addr = IBuf_state;
  assign IBuf_cov_write_mask = 1'h1;
  assign IBuf_cov_write_en = 1'h1;
  assign nBufValid_shl = nBufValid;
  assign nBufValid_pad = {1'h0,nBufValid_shl};
  assign buf__replay_shl = {buf__replay, 1'h0};
  assign buf__replay_pad = buf__replay_shl;
  assign IBuf_xor0 = nBufValid_pad ^ buf__replay_pad;
  assign RVCExpander_sum = IBuf_covSum + RVCExpander_io_covSum;
  assign io_covSum = RVCExpander_sum;
  assign stopEn0 = ~_T_112;
  assign RVCExpander_metaAssert_wire = RVCExpander_metaAssert;
  assign IBuf_or0 = stopEn0 | RVCExpander_metaAssert_wire;
  assign metaAssert = IBuf_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  nBufValid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  buf__pc = _RAND_1[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  buf__data = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  buf__xcpt_pf_inst = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  buf__xcpt_ae_inst = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  buf__replay = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  ibufBTBResp_entry = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ibufBTBResp_bht_history = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  IBuf_state = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    IBuf_cov[initvar] = _RAND_9[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  IBuf_covSum = _RAND_10[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  IBuf_metaAssert = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      nBufValid <= 1'h0;
    end else if (reset) begin
      nBufValid <= 1'h0;
    end else begin
      nBufValid <= _GEN_46[0];
    end
    if (metaReset) begin
      buf__pc <= 40'h0;
    end else if (io_inst_0_ready) begin
      if (_T_55) begin
        buf__pc <= _T_73;
      end
    end
    if (metaReset) begin
      buf__data <= 32'h0;
    end else if (io_inst_0_ready) begin
      if (_T_55) begin
        buf__data <= {{16'd0}, _T_65[15:0]};
      end
    end
    if (metaReset) begin
      buf__xcpt_pf_inst <= 1'h0;
    end else if (io_inst_0_ready) begin
      if (_T_55) begin
        buf__xcpt_pf_inst <= io_imem_bits_xcpt_pf_inst;
      end
    end
    if (metaReset) begin
      buf__xcpt_ae_inst <= 1'h0;
    end else if (io_inst_0_ready) begin
      if (_T_55) begin
        buf__xcpt_ae_inst <= io_imem_bits_xcpt_ae_inst;
      end
    end
    if (metaReset) begin
      buf__replay <= 1'h0;
    end else if (io_inst_0_ready) begin
      if (_T_55) begin
        buf__replay <= io_imem_bits_replay;
      end
    end
    if (metaReset) begin
      ibufBTBResp_entry <= 5'h0;
    end else if (io_inst_0_ready) begin
      if (_T_55) begin
        ibufBTBResp_entry <= io_imem_bits_btb_entry;
      end
    end
    if (metaReset) begin
      ibufBTBResp_bht_history <= 8'h0;
    end else if (io_inst_0_ready) begin
      if (_T_55) begin
        ibufBTBResp_bht_history <= io_imem_bits_btb_bht_history;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_112) begin
          $fwrite(32'h80000002,"Assertion failed\n    at IBuf.scala:79 assert(!io.imem.valid || !io.imem.bits.btb.taken || io.imem.bits.btb.bridx >= pcWordBits)\n"); // @[IBuf.scala 79:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_112) begin
          $fatal; // @[IBuf.scala 79:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    IBuf_state <= IBuf_xor0;
    if (!(IBuf_cov_read_data)) begin
      IBuf_covSum <= IBuf_covSum + 1'h1;
    end
    if (metaReset) begin
      IBuf_metaAssert <= 1'h0;
    end else begin
      IBuf_metaAssert <= IBuf_metaAssert | IBuf_or0;
    end
  end
  always @(posedge clock) begin
    if(IBuf_cov_write_en & IBuf_cov_write_mask) begin
      IBuf_cov[IBuf_cov_write_addr] <= IBuf_cov_write_data; // @[Coverage map for IBuf]
    end
  end
endmodule
module CSRFile(
  input         clock,
  input         reset,
  input         io_ungated_clock,
  input         io_interrupts_debug,
  input         io_interrupts_mtip,
  input         io_interrupts_msip,
  input         io_interrupts_meip,
  input         io_interrupts_seip,
  input  [1:0]  io_hartid,
  input  [11:0] io_rw_addr,
  input  [2:0]  io_rw_cmd,
  output [63:0] io_rw_rdata,
  input  [63:0] io_rw_wdata,
  output        io_pcode_req_valid,
  output [1:0]  io_pcode_req_bits_id,
  output [19:0] io_pcode_req_bits_value_base,
  output [9:0]  io_pcode_req_bits_value_mask,
  output        io_pcode_req_bits_value_valid,
  output        io_pcode_req_bits_value_locked,
  output [26:0] io_vpoffset_req_bits_value,
  input  [11:0] io_decode_0_csr,
  output        io_decode_0_fp_illegal,
  output        io_decode_0_fp_csr,
  output        io_decode_0_read_illegal,
  output        io_decode_0_write_illegal,
  output        io_decode_0_write_flush,
  output        io_decode_0_system_illegal,
  output        io_csr_stall,
  output        io_eret,
  output        io_singleStep,
  output        io_status_debug,
  output [31:0] io_status_isa,
  output [1:0]  io_status_dprv,
  output [1:0]  io_status_prv,
  output        io_status_sd,
  output [26:0] io_status_zero2,
  output [1:0]  io_status_sxl,
  output [1:0]  io_status_uxl,
  output        io_status_sd_rv32,
  output [7:0]  io_status_zero1,
  output        io_status_tsr,
  output        io_status_tw,
  output        io_status_tvm,
  output        io_status_mxr,
  output        io_status_sum,
  output        io_status_mprv,
  output [1:0]  io_status_xs,
  output [1:0]  io_status_fs,
  output [1:0]  io_status_mpp,
  output [1:0]  io_status_hpp,
  output        io_status_spp,
  output        io_status_mpie,
  output        io_status_hpie,
  output        io_status_spie,
  output        io_status_upie,
  output        io_status_mie,
  output        io_status_hie,
  output        io_status_sie,
  output        io_status_uie,
  output [3:0]  io_ptbr_mode,
  output [43:0] io_ptbr_ppn,
  output [39:0] io_evec,
  input         io_exception,
  input         io_retire,
  input  [63:0] io_cause,
  input  [39:0] io_pc,
  input  [39:0] io_tval,
  output [2:0]  io_fcsr_rm,
  input         io_fcsr_flags_valid,
  input  [4:0]  io_fcsr_flags_bits,
  output        io_interrupt,
  output [63:0] io_interrupt_cause,
  output        io_bp_0_control_action,
  output [1:0]  io_bp_0_control_tmatch,
  output        io_bp_0_control_m,
  output        io_bp_0_control_s,
  output        io_bp_0_control_u,
  output        io_bp_0_control_x,
  output        io_bp_0_control_w,
  output        io_bp_0_control_r,
  output [38:0] io_bp_0_address,
  output        io_pmp_0_cfg_l,
  output [1:0]  io_pmp_0_cfg_a,
  output        io_pmp_0_cfg_x,
  output        io_pmp_0_cfg_w,
  output        io_pmp_0_cfg_r,
  output [29:0] io_pmp_0_addr,
  output [31:0] io_pmp_0_mask,
  output        io_pmp_1_cfg_l,
  output [1:0]  io_pmp_1_cfg_a,
  output        io_pmp_1_cfg_x,
  output        io_pmp_1_cfg_w,
  output        io_pmp_1_cfg_r,
  output [29:0] io_pmp_1_addr,
  output [31:0] io_pmp_1_mask,
  output        io_pmp_2_cfg_l,
  output [1:0]  io_pmp_2_cfg_a,
  output        io_pmp_2_cfg_x,
  output        io_pmp_2_cfg_w,
  output        io_pmp_2_cfg_r,
  output [29:0] io_pmp_2_addr,
  output [31:0] io_pmp_2_mask,
  output        io_pmp_3_cfg_l,
  output [1:0]  io_pmp_3_cfg_a,
  output        io_pmp_3_cfg_x,
  output        io_pmp_3_cfg_w,
  output        io_pmp_3_cfg_r,
  output [29:0] io_pmp_3_addr,
  output [31:0] io_pmp_3_mask,
  output        io_pmp_4_cfg_l,
  output [1:0]  io_pmp_4_cfg_a,
  output        io_pmp_4_cfg_x,
  output        io_pmp_4_cfg_w,
  output        io_pmp_4_cfg_r,
  output [29:0] io_pmp_4_addr,
  output [31:0] io_pmp_4_mask,
  output        io_pmp_5_cfg_l,
  output [1:0]  io_pmp_5_cfg_a,
  output        io_pmp_5_cfg_x,
  output        io_pmp_5_cfg_w,
  output        io_pmp_5_cfg_r,
  output [29:0] io_pmp_5_addr,
  output [31:0] io_pmp_5_mask,
  output        io_pmp_6_cfg_l,
  output [1:0]  io_pmp_6_cfg_a,
  output        io_pmp_6_cfg_x,
  output        io_pmp_6_cfg_w,
  output        io_pmp_6_cfg_r,
  output [29:0] io_pmp_6_addr,
  output [31:0] io_pmp_6_mask,
  output        io_pmp_7_cfg_l,
  output [1:0]  io_pmp_7_cfg_a,
  output        io_pmp_7_cfg_x,
  output        io_pmp_7_cfg_w,
  output        io_pmp_7_cfg_r,
  output [29:0] io_pmp_7_addr,
  output [31:0] io_pmp_7_mask,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [1:0] reg_mstatus_prv; // @[CSR.scala 272:24]
  reg [31:0] _RAND_0;
  reg  reg_mstatus_tsr; // @[CSR.scala 272:24]
  reg [31:0] _RAND_1;
  reg  reg_mstatus_tw; // @[CSR.scala 272:24]
  reg [31:0] _RAND_2;
  reg  reg_mstatus_tvm; // @[CSR.scala 272:24]
  reg [31:0] _RAND_3;
  reg  reg_mstatus_mxr; // @[CSR.scala 272:24]
  reg [31:0] _RAND_4;
  reg  reg_mstatus_sum; // @[CSR.scala 272:24]
  reg [31:0] _RAND_5;
  reg  reg_mstatus_mprv; // @[CSR.scala 272:24]
  reg [31:0] _RAND_6;
  reg [1:0] reg_mstatus_fs; // @[CSR.scala 272:24]
  reg [31:0] _RAND_7;
  reg [1:0] reg_mstatus_mpp; // @[CSR.scala 272:24]
  reg [31:0] _RAND_8;
  reg  reg_mstatus_spp; // @[CSR.scala 272:24]
  reg [31:0] _RAND_9;
  reg  reg_mstatus_mpie; // @[CSR.scala 272:24]
  reg [31:0] _RAND_10;
  reg  reg_mstatus_spie; // @[CSR.scala 272:24]
  reg [31:0] _RAND_11;
  reg  reg_mstatus_mie; // @[CSR.scala 272:24]
  reg [31:0] _RAND_12;
  reg  reg_mstatus_sie; // @[CSR.scala 272:24]
  reg [31:0] _RAND_13;
  wire  system_insn; // @[CSR.scala 581:31]
  wire [31:0] _T_1137; // @[CSR.scala 590:92]
  wire [31:0] _T_1144; // @[Decode.scala 14:65]
  wire  _T_1145; // @[Decode.scala 14:121]
  wire [31:0] _T_1146; // @[Decode.scala 14:65]
  wire  _T_1147; // @[Decode.scala 14:121]
  wire  _T_1149; // @[Decode.scala 15:30]
  wire  insn_ret; // @[CSR.scala 590:159]
  reg [1:0] reg_dcsr_prv; // @[CSR.scala 280:21]
  reg [31:0] _RAND_14;
  wire [1:0] _GEN_125; // @[CSR.scala 725:53]
  wire [1:0] _GEN_134; // @[CSR.scala 719:44]
  wire [31:0] _T_1138; // @[Decode.scala 14:65]
  wire  _T_1139; // @[Decode.scala 14:121]
  wire  insn_call; // @[CSR.scala 590:159]
  wire  _T_1142; // @[Decode.scala 14:121]
  wire  insn_break; // @[CSR.scala 590:159]
  wire  _T_1627; // @[CSR.scala 655:29]
  wire  exception; // @[CSR.scala 655:43]
  reg  reg_singleStepped; // @[CSR.scala 324:30]
  reg [31:0] _RAND_15;
  wire [3:0] _GEN_727; // @[CSR.scala 619:36]
  wire [3:0] _T_1572; // @[CSR.scala 619:36]
  wire [63:0] _T_1573; // @[CSR.scala 620:14]
  wire [63:0] cause; // @[CSR.scala 619:8]
  wire [7:0] cause_lsbs; // @[CSR.scala 621:25]
  wire  _T_1575; // @[CSR.scala 622:53]
  wire  causeIsDebugInt; // @[CSR.scala 622:39]
  wire  _T_1587; // @[CSR.scala 625:60]
  wire  causeIsDebugTrigger; // @[CSR.scala 623:44]
  wire  _T_1588; // @[CSR.scala 625:79]
  wire  _T_1581; // @[CSR.scala 624:42]
  reg  reg_dcsr_ebreakm; // @[CSR.scala 280:21]
  reg [31:0] _RAND_16;
  reg  reg_dcsr_ebreaks; // @[CSR.scala 280:21]
  reg [31:0] _RAND_17;
  reg  reg_dcsr_ebreaku; // @[CSR.scala 280:21]
  reg [31:0] _RAND_18;
  wire [3:0] _T_1584; // @[Cat.scala 30:58]
  wire [3:0] _T_1585; // @[CSR.scala 624:134]
  wire  causeIsDebugBreak; // @[CSR.scala 624:56]
  wire  _T_1589; // @[CSR.scala 625:102]
  reg  reg_debug; // @[CSR.scala 321:22]
  reg [31:0] _RAND_19;
  wire  trapToDebug; // @[CSR.scala 625:123]
  wire [1:0] _GEN_74; // @[CSR.scala 672:25]
  wire  _T_1592; // @[CSR.scala 627:51]
  reg [63:0] reg_mideleg; // @[CSR.scala 331:24]
  reg [63:0] _RAND_20;
  wire [63:0] _T_1595; // @[CSR.scala 627:93]
  reg [63:0] reg_medeleg; // @[CSR.scala 332:24]
  reg [63:0] _RAND_21;
  wire [63:0] _T_1597; // @[CSR.scala 627:118]
  wire  _T_1599; // @[CSR.scala 627:66]
  wire  delegate; // @[CSR.scala 627:60]
  wire [1:0] _GEN_82; // @[CSR.scala 679:27]
  wire [1:0] _GEN_93; // @[CSR.scala 671:24]
  wire [1:0] _GEN_111; // @[CSR.scala 670:20]
  wire [1:0] new_prv; // @[CSR.scala 718:19]
  wire  _T_172; // @[CSR.scala 1035:27]
  reg [2:0] reg_dcsr_cause; // @[CSR.scala 280:21]
  reg [31:0] _RAND_22;
  reg  reg_dcsr_step; // @[CSR.scala 280:21]
  reg [31:0] _RAND_23;
  reg [39:0] reg_dpc; // @[CSR.scala 322:20]
  reg [63:0] _RAND_24;
  reg [63:0] reg_dscratch; // @[CSR.scala 323:25]
  reg [63:0] _RAND_25;
  reg  reg_bp_0_control_dmode; // @[CSR.scala 327:19]
  reg [31:0] _RAND_26;
  reg  reg_bp_0_control_action; // @[CSR.scala 327:19]
  reg [31:0] _RAND_27;
  reg [1:0] reg_bp_0_control_tmatch; // @[CSR.scala 327:19]
  reg [31:0] _RAND_28;
  reg  reg_bp_0_control_m; // @[CSR.scala 327:19]
  reg [31:0] _RAND_29;
  reg  reg_bp_0_control_s; // @[CSR.scala 327:19]
  reg [31:0] _RAND_30;
  reg  reg_bp_0_control_u; // @[CSR.scala 327:19]
  reg [31:0] _RAND_31;
  reg  reg_bp_0_control_x; // @[CSR.scala 327:19]
  reg [31:0] _RAND_32;
  reg  reg_bp_0_control_w; // @[CSR.scala 327:19]
  reg [31:0] _RAND_33;
  reg  reg_bp_0_control_r; // @[CSR.scala 327:19]
  reg [31:0] _RAND_34;
  reg [38:0] reg_bp_0_address; // @[CSR.scala 327:19]
  reg [63:0] _RAND_35;
  reg  reg_pmp_0_cfg_l; // @[CSR.scala 328:20]
  reg [31:0] _RAND_36;
  reg [1:0] reg_pmp_0_cfg_a; // @[CSR.scala 328:20]
  reg [31:0] _RAND_37;
  reg  reg_pmp_0_cfg_x; // @[CSR.scala 328:20]
  reg [31:0] _RAND_38;
  reg  reg_pmp_0_cfg_w; // @[CSR.scala 328:20]
  reg [31:0] _RAND_39;
  reg  reg_pmp_0_cfg_r; // @[CSR.scala 328:20]
  reg [31:0] _RAND_40;
  reg [29:0] reg_pmp_0_addr; // @[CSR.scala 328:20]
  reg [31:0] _RAND_41;
  reg  reg_pmp_1_cfg_l; // @[CSR.scala 328:20]
  reg [31:0] _RAND_42;
  reg [1:0] reg_pmp_1_cfg_a; // @[CSR.scala 328:20]
  reg [31:0] _RAND_43;
  reg  reg_pmp_1_cfg_x; // @[CSR.scala 328:20]
  reg [31:0] _RAND_44;
  reg  reg_pmp_1_cfg_w; // @[CSR.scala 328:20]
  reg [31:0] _RAND_45;
  reg  reg_pmp_1_cfg_r; // @[CSR.scala 328:20]
  reg [31:0] _RAND_46;
  reg [29:0] reg_pmp_1_addr; // @[CSR.scala 328:20]
  reg [31:0] _RAND_47;
  reg  reg_pmp_2_cfg_l; // @[CSR.scala 328:20]
  reg [31:0] _RAND_48;
  reg [1:0] reg_pmp_2_cfg_a; // @[CSR.scala 328:20]
  reg [31:0] _RAND_49;
  reg  reg_pmp_2_cfg_x; // @[CSR.scala 328:20]
  reg [31:0] _RAND_50;
  reg  reg_pmp_2_cfg_w; // @[CSR.scala 328:20]
  reg [31:0] _RAND_51;
  reg  reg_pmp_2_cfg_r; // @[CSR.scala 328:20]
  reg [31:0] _RAND_52;
  reg [29:0] reg_pmp_2_addr; // @[CSR.scala 328:20]
  reg [31:0] _RAND_53;
  reg  reg_pmp_3_cfg_l; // @[CSR.scala 328:20]
  reg [31:0] _RAND_54;
  reg [1:0] reg_pmp_3_cfg_a; // @[CSR.scala 328:20]
  reg [31:0] _RAND_55;
  reg  reg_pmp_3_cfg_x; // @[CSR.scala 328:20]
  reg [31:0] _RAND_56;
  reg  reg_pmp_3_cfg_w; // @[CSR.scala 328:20]
  reg [31:0] _RAND_57;
  reg  reg_pmp_3_cfg_r; // @[CSR.scala 328:20]
  reg [31:0] _RAND_58;
  reg [29:0] reg_pmp_3_addr; // @[CSR.scala 328:20]
  reg [31:0] _RAND_59;
  reg  reg_pmp_4_cfg_l; // @[CSR.scala 328:20]
  reg [31:0] _RAND_60;
  reg [1:0] reg_pmp_4_cfg_a; // @[CSR.scala 328:20]
  reg [31:0] _RAND_61;
  reg  reg_pmp_4_cfg_x; // @[CSR.scala 328:20]
  reg [31:0] _RAND_62;
  reg  reg_pmp_4_cfg_w; // @[CSR.scala 328:20]
  reg [31:0] _RAND_63;
  reg  reg_pmp_4_cfg_r; // @[CSR.scala 328:20]
  reg [31:0] _RAND_64;
  reg [29:0] reg_pmp_4_addr; // @[CSR.scala 328:20]
  reg [31:0] _RAND_65;
  reg  reg_pmp_5_cfg_l; // @[CSR.scala 328:20]
  reg [31:0] _RAND_66;
  reg [1:0] reg_pmp_5_cfg_a; // @[CSR.scala 328:20]
  reg [31:0] _RAND_67;
  reg  reg_pmp_5_cfg_x; // @[CSR.scala 328:20]
  reg [31:0] _RAND_68;
  reg  reg_pmp_5_cfg_w; // @[CSR.scala 328:20]
  reg [31:0] _RAND_69;
  reg  reg_pmp_5_cfg_r; // @[CSR.scala 328:20]
  reg [31:0] _RAND_70;
  reg [29:0] reg_pmp_5_addr; // @[CSR.scala 328:20]
  reg [31:0] _RAND_71;
  reg  reg_pmp_6_cfg_l; // @[CSR.scala 328:20]
  reg [31:0] _RAND_72;
  reg [1:0] reg_pmp_6_cfg_a; // @[CSR.scala 328:20]
  reg [31:0] _RAND_73;
  reg  reg_pmp_6_cfg_x; // @[CSR.scala 328:20]
  reg [31:0] _RAND_74;
  reg  reg_pmp_6_cfg_w; // @[CSR.scala 328:20]
  reg [31:0] _RAND_75;
  reg  reg_pmp_6_cfg_r; // @[CSR.scala 328:20]
  reg [31:0] _RAND_76;
  reg [29:0] reg_pmp_6_addr; // @[CSR.scala 328:20]
  reg [31:0] _RAND_77;
  reg  reg_pmp_7_cfg_l; // @[CSR.scala 328:20]
  reg [31:0] _RAND_78;
  reg [1:0] reg_pmp_7_cfg_a; // @[CSR.scala 328:20]
  reg [31:0] _RAND_79;
  reg  reg_pmp_7_cfg_x; // @[CSR.scala 328:20]
  reg [31:0] _RAND_80;
  reg  reg_pmp_7_cfg_w; // @[CSR.scala 328:20]
  reg [31:0] _RAND_81;
  reg  reg_pmp_7_cfg_r; // @[CSR.scala 328:20]
  reg [31:0] _RAND_82;
  reg [29:0] reg_pmp_7_addr; // @[CSR.scala 328:20]
  reg [31:0] _RAND_83;
  reg [63:0] reg_mie; // @[CSR.scala 330:20]
  reg [63:0] _RAND_84;
  reg  reg_mip_seip; // @[CSR.scala 333:20]
  reg [31:0] _RAND_85;
  reg  reg_mip_stip; // @[CSR.scala 333:20]
  reg [31:0] _RAND_86;
  reg  reg_mip_ssip; // @[CSR.scala 333:20]
  reg [31:0] _RAND_87;
  reg [39:0] reg_mepc; // @[CSR.scala 334:21]
  reg [63:0] _RAND_88;
  reg [63:0] reg_mcause; // @[CSR.scala 335:23]
  reg [63:0] _RAND_89;
  reg [39:0] reg_mbadaddr; // @[CSR.scala 336:25]
  reg [63:0] _RAND_90;
  reg [63:0] reg_mscratch; // @[CSR.scala 337:25]
  reg [63:0] _RAND_91;
  reg [31:0] reg_mtvec; // @[CSR.scala 340:27]
  reg [31:0] _RAND_92;
  reg [31:0] reg_mcounteren; // @[CSR.scala 343:27]
  reg [31:0] _RAND_93;
  reg [31:0] reg_scounteren; // @[CSR.scala 344:27]
  reg [31:0] _RAND_94;
  reg [39:0] reg_sepc; // @[CSR.scala 347:21]
  reg [63:0] _RAND_95;
  reg [63:0] reg_scause; // @[CSR.scala 348:23]
  reg [63:0] _RAND_96;
  reg [39:0] reg_sbadaddr; // @[CSR.scala 349:25]
  reg [63:0] _RAND_97;
  reg [63:0] reg_sscratch; // @[CSR.scala 350:25]
  reg [63:0] _RAND_98;
  reg [38:0] reg_stvec; // @[CSR.scala 351:22]
  reg [63:0] _RAND_99;
  reg [3:0] reg_sptbr_mode; // @[CSR.scala 352:22]
  reg [31:0] _RAND_100;
  reg [43:0] reg_sptbr_ppn; // @[CSR.scala 352:22]
  reg [63:0] _RAND_101;
  reg  reg_wfi; // @[CSR.scala 353:50]
  reg [31:0] _RAND_102;
  reg [4:0] reg_fflags; // @[CSR.scala 355:23]
  reg [31:0] _RAND_103;
  reg [2:0] reg_frm; // @[CSR.scala 356:20]
  reg [31:0] _RAND_104;
  reg [5:0] _T_286; // @[Counters.scala 46:37]
  reg [31:0] _RAND_105;
  wire [5:0] _GEN_728; // @[Counters.scala 47:33]
  wire [6:0] _T_287; // @[Counters.scala 47:33]
  reg [57:0] _T_289; // @[Counters.scala 51:27]
  reg [63:0] _RAND_106;
  wire [57:0] _T_292; // @[Counters.scala 52:43]
  wire [63:0] _T_293; // @[Cat.scala 30:58]
  reg [5:0] _T_296; // @[Counters.scala 46:37]
  reg [31:0] _RAND_107;
  wire [5:0] _GEN_729; // @[Counters.scala 47:33]
  wire [6:0] _T_297; // @[Counters.scala 47:33]
  reg [57:0] _T_299; // @[Counters.scala 51:27]
  reg [63:0] _RAND_108;
  wire [57:0] _T_302; // @[Counters.scala 52:43]
  wire [63:0] _T_303; // @[Cat.scala 30:58]
  reg  _T_310; // @[CSR.scala 370:67]
  reg [31:0] _RAND_109;
  wire  mip_seip; // @[CSR.scala 370:57]
  wire [7:0] _T_318; // @[CSR.scala 372:22]
  wire [15:0] _T_326; // @[CSR.scala 372:22]
  wire [15:0] read_mip; // @[CSR.scala 372:29]
  wire [63:0] _GEN_730; // @[CSR.scala 375:56]
  wire [63:0] pending_interrupts; // @[CSR.scala 375:56]
  wire [14:0] d_interrupts; // @[CSR.scala 376:42]
  wire  _T_329; // @[CSR.scala 377:51]
  wire [63:0] _T_331; // @[CSR.scala 377:93]
  wire [63:0] m_interrupts; // @[CSR.scala 377:25]
  wire  _T_333; // @[CSR.scala 378:42]
  wire  _T_334; // @[CSR.scala 378:70]
  wire  _T_335; // @[CSR.scala 378:80]
  wire  _T_336; // @[CSR.scala 378:50]
  wire [63:0] _T_337; // @[CSR.scala 378:120]
  wire [63:0] s_interrupts; // @[CSR.scala 378:25]
  wire  _T_376; // @[CSR.scala 1025:90]
  wire  _T_377; // @[CSR.scala 1025:90]
  wire  _T_378; // @[CSR.scala 1025:90]
  wire  _T_379; // @[CSR.scala 1025:90]
  wire  _T_380; // @[CSR.scala 1025:90]
  wire  _T_381; // @[CSR.scala 1025:90]
  wire  _T_382; // @[CSR.scala 1025:90]
  wire  _T_383; // @[CSR.scala 1025:90]
  wire  _T_384; // @[CSR.scala 1025:90]
  wire  _T_385; // @[CSR.scala 1025:90]
  wire  _T_386; // @[CSR.scala 1025:90]
  wire  _T_387; // @[CSR.scala 1025:90]
  wire  _T_388; // @[CSR.scala 1025:90]
  wire  _T_389; // @[CSR.scala 1025:90]
  wire  _T_390; // @[CSR.scala 1025:90]
  wire  _T_391; // @[CSR.scala 1025:90]
  wire  _T_392; // @[CSR.scala 1025:90]
  wire  _T_393; // @[CSR.scala 1025:90]
  wire  _T_394; // @[CSR.scala 1025:90]
  wire  _T_395; // @[CSR.scala 1025:90]
  wire  _T_396; // @[CSR.scala 1025:90]
  wire  _T_397; // @[CSR.scala 1025:90]
  wire  _T_398; // @[CSR.scala 1025:90]
  wire  _T_399; // @[CSR.scala 1025:90]
  wire  _T_400; // @[CSR.scala 1025:90]
  wire  _T_401; // @[CSR.scala 1025:90]
  wire  _T_402; // @[CSR.scala 1025:90]
  wire  _T_403; // @[CSR.scala 1025:90]
  wire  _T_404; // @[CSR.scala 1025:90]
  wire  _T_405; // @[CSR.scala 1025:90]
  wire  _T_406; // @[CSR.scala 1025:90]
  wire  _T_407; // @[CSR.scala 1025:90]
  wire  _T_408; // @[CSR.scala 1025:90]
  wire  _T_409; // @[CSR.scala 1025:90]
  wire  _T_410; // @[CSR.scala 1025:90]
  wire  _T_411; // @[CSR.scala 1025:90]
  wire  anyInterrupt; // @[CSR.scala 1025:90]
  wire [2:0] _T_450; // @[Mux.scala 31:69]
  wire [3:0] _T_451; // @[Mux.scala 31:69]
  wire [3:0] _T_452; // @[Mux.scala 31:69]
  wire [3:0] _T_453; // @[Mux.scala 31:69]
  wire [3:0] _T_454; // @[Mux.scala 31:69]
  wire [3:0] _T_455; // @[Mux.scala 31:69]
  wire [3:0] _T_456; // @[Mux.scala 31:69]
  wire [3:0] _T_457; // @[Mux.scala 31:69]
  wire [3:0] _T_458; // @[Mux.scala 31:69]
  wire [3:0] _T_459; // @[Mux.scala 31:69]
  wire [3:0] _T_460; // @[Mux.scala 31:69]
  wire [3:0] _T_461; // @[Mux.scala 31:69]
  wire [3:0] _T_462; // @[Mux.scala 31:69]
  wire [3:0] _T_463; // @[Mux.scala 31:69]
  wire [3:0] _T_464; // @[Mux.scala 31:69]
  wire [3:0] _T_465; // @[Mux.scala 31:69]
  wire [3:0] _T_466; // @[Mux.scala 31:69]
  wire [3:0] _T_467; // @[Mux.scala 31:69]
  wire [3:0] _T_468; // @[Mux.scala 31:69]
  wire [3:0] _T_469; // @[Mux.scala 31:69]
  wire [3:0] _T_470; // @[Mux.scala 31:69]
  wire [3:0] _T_471; // @[Mux.scala 31:69]
  wire [3:0] _T_472; // @[Mux.scala 31:69]
  wire [3:0] _T_473; // @[Mux.scala 31:69]
  wire [3:0] _T_474; // @[Mux.scala 31:69]
  wire [3:0] _T_475; // @[Mux.scala 31:69]
  wire [3:0] _T_476; // @[Mux.scala 31:69]
  wire [3:0] _T_477; // @[Mux.scala 31:69]
  wire [3:0] _T_478; // @[Mux.scala 31:69]
  wire [3:0] _T_479; // @[Mux.scala 31:69]
  wire [3:0] _T_480; // @[Mux.scala 31:69]
  wire [3:0] _T_481; // @[Mux.scala 31:69]
  wire [3:0] _T_482; // @[Mux.scala 31:69]
  wire [3:0] _T_483; // @[Mux.scala 31:69]
  wire [3:0] _T_484; // @[Mux.scala 31:69]
  wire [3:0] _T_485; // @[Mux.scala 31:69]
  wire [3:0] whichInterrupt; // @[Mux.scala 31:69]
  wire [63:0] _GEN_731; // @[CSR.scala 381:43]
  wire  _T_488; // @[CSR.scala 382:33]
  wire  _T_489; // @[CSR.scala 382:51]
  wire [30:0] _T_495; // @[Cat.scala 30:58]
  wire [30:0] _T_498; // @[PMP.scala 52:23]
  wire [30:0] _T_500; // @[PMP.scala 52:14]
  wire [32:0] _T_501; // @[Cat.scala 30:58]
  wire [30:0] _T_505; // @[Cat.scala 30:58]
  wire [30:0] _T_508; // @[PMP.scala 52:23]
  wire [30:0] _T_510; // @[PMP.scala 52:14]
  wire [32:0] _T_511; // @[Cat.scala 30:58]
  wire [30:0] _T_515; // @[Cat.scala 30:58]
  wire [30:0] _T_518; // @[PMP.scala 52:23]
  wire [30:0] _T_520; // @[PMP.scala 52:14]
  wire [32:0] _T_521; // @[Cat.scala 30:58]
  wire [30:0] _T_525; // @[Cat.scala 30:58]
  wire [30:0] _T_528; // @[PMP.scala 52:23]
  wire [30:0] _T_530; // @[PMP.scala 52:14]
  wire [32:0] _T_531; // @[Cat.scala 30:58]
  wire [30:0] _T_535; // @[Cat.scala 30:58]
  wire [30:0] _T_538; // @[PMP.scala 52:23]
  wire [30:0] _T_540; // @[PMP.scala 52:14]
  wire [32:0] _T_541; // @[Cat.scala 30:58]
  wire [30:0] _T_545; // @[Cat.scala 30:58]
  wire [30:0] _T_548; // @[PMP.scala 52:23]
  wire [30:0] _T_550; // @[PMP.scala 52:14]
  wire [32:0] _T_551; // @[Cat.scala 30:58]
  wire [30:0] _T_555; // @[Cat.scala 30:58]
  wire [30:0] _T_558; // @[PMP.scala 52:23]
  wire [30:0] _T_560; // @[PMP.scala 52:14]
  wire [32:0] _T_561; // @[Cat.scala 30:58]
  wire [30:0] _T_565; // @[Cat.scala 30:58]
  wire [30:0] _T_568; // @[PMP.scala 52:23]
  wire [30:0] _T_570; // @[PMP.scala 52:14]
  wire [32:0] _T_571; // @[Cat.scala 30:58]
  reg [63:0] reg_misa; // @[CSR.scala 398:21]
  reg [63:0] _RAND_110;
  wire [6:0] _T_578; // @[CSR.scala 399:38]
  wire [17:0] _T_585; // @[CSR.scala 399:38]
  wire [13:0] _T_591; // @[CSR.scala 399:38]
  wire [100:0] _T_600; // @[CSR.scala 399:38]
  wire [63:0] read_mstatus; // @[CSR.scala 399:40]
  wire [6:0] _T_607; // @[CSR.scala 403:48]
  wire [63:0] _T_615; // @[CSR.scala 403:48]
  wire [24:0] _T_619; // @[Bitwise.scala 72:12]
  wire [63:0] _T_620; // @[Cat.scala 30:58]
  wire [1:0] _T_623; // @[CSR.scala 1053:36]
  wire [39:0] _GEN_732; // @[CSR.scala 1053:31]
  wire [39:0] _T_624; // @[CSR.scala 1053:31]
  wire  _T_626; // @[package.scala 106:38]
  wire [23:0] _T_628; // @[Bitwise.scala 72:12]
  wire [63:0] _T_629; // @[Cat.scala 30:58]
  wire [23:0] _T_632; // @[Bitwise.scala 72:12]
  wire [63:0] _T_633; // @[Cat.scala 30:58]
  wire [11:0] _T_639; // @[CSR.scala 417:27]
  wire [31:0] _T_646; // @[CSR.scala 417:27]
  wire [39:0] _T_650; // @[CSR.scala 1053:31]
  wire  _T_652; // @[package.scala 106:38]
  wire [23:0] _T_654; // @[Bitwise.scala 72:12]
  wire [63:0] _T_655; // @[Cat.scala 30:58]
  wire [7:0] _T_656; // @[Cat.scala 30:58]
  reg [26:0] vpoffset_reg; // @[CSR.scala 470:25]
  reg [31:0] _RAND_111;
  reg  pcode_regs_0_locked; // @[CSR.scala 473:23]
  reg [31:0] _RAND_112;
  reg  pcode_regs_1_locked; // @[CSR.scala 473:23]
  reg [31:0] _RAND_113;
  reg  pcode_regs_2_locked; // @[CSR.scala 473:23]
  reg [31:0] _RAND_114;
  reg  pcode_regs_3_locked; // @[CSR.scala 473:23]
  reg [31:0] _RAND_115;
  reg  pcode_update_valid; // @[CSR.scala 487:25]
  reg [31:0] _RAND_116;
  reg [1:0] pcode_update_bits_id; // @[CSR.scala 487:25]
  reg [31:0] _RAND_117;
  reg [19:0] pcode_update_bits_value_base; // @[CSR.scala 487:25]
  reg [31:0] _RAND_118;
  reg [9:0] pcode_update_bits_value_mask; // @[CSR.scala 487:25]
  reg [31:0] _RAND_119;
  reg  pcode_update_bits_value_valid; // @[CSR.scala 487:25]
  reg [31:0] _RAND_120;
  reg  pcode_update_bits_value_locked; // @[CSR.scala 487:25]
  reg [31:0] _RAND_121;
  reg [26:0] vpoffset_update_bits_value; // @[CSR.scala 490:28]
  reg [31:0] _RAND_122;
  wire [31:0] _T_771; // @[Cat.scala 30:58]
  wire [31:0] _T_774; // @[Cat.scala 30:58]
  wire [31:0] _T_777; // @[Cat.scala 30:58]
  wire [31:0] _T_780; // @[Cat.scala 30:58]
  wire [63:0] _T_781; // @[CSR.scala 527:28]
  wire [63:0] _T_782; // @[CSR.scala 528:29]
  wire [6:0] _T_824; // @[CSR.scala 541:57]
  wire [17:0] _T_831; // @[CSR.scala 541:57]
  wire [13:0] _T_837; // @[CSR.scala 541:57]
  wire [100:0] _T_846; // @[CSR.scala 541:57]
  wire [23:0] _T_850; // @[Bitwise.scala 72:12]
  wire [63:0] _T_851; // @[Cat.scala 30:58]
  wire [63:0] _T_853; // @[CSR.scala 547:45]
  wire [39:0] _T_857; // @[CSR.scala 1053:31]
  wire  _T_859; // @[package.scala 106:38]
  wire [23:0] _T_861; // @[Bitwise.scala 72:12]
  wire [63:0] _T_862; // @[Cat.scala 30:58]
  wire [24:0] _T_865; // @[Bitwise.scala 72:12]
  wire [63:0] _T_866; // @[Cat.scala 30:58]
  wire [7:0] _T_885; // @[package.scala 35:38]
  wire [7:0] _T_895; // @[package.scala 35:38]
  wire [7:0] _T_905; // @[package.scala 35:38]
  wire [7:0] _T_915; // @[package.scala 35:38]
  wire [15:0] _T_921; // @[Cat.scala 30:58]
  wire [31:0] _T_923; // @[Cat.scala 30:58]
  wire [15:0] _T_924; // @[Cat.scala 30:58]
  wire [63:0] _T_927; // @[Cat.scala 30:58]
  wire  _T_980; // @[CSR.scala 578:73]
  wire  _T_981; // @[CSR.scala 578:73]
  wire  _T_982; // @[CSR.scala 578:73]
  wire  _T_983; // @[CSR.scala 578:73]
  wire  _T_984; // @[CSR.scala 578:73]
  wire  _T_985; // @[CSR.scala 578:73]
  wire  _T_986; // @[CSR.scala 578:73]
  wire  _T_987; // @[CSR.scala 578:73]
  wire  _T_988; // @[CSR.scala 578:73]
  wire  _T_989; // @[CSR.scala 578:73]
  wire  _T_990; // @[CSR.scala 578:73]
  wire  _T_991; // @[CSR.scala 578:73]
  wire  _T_992; // @[CSR.scala 578:73]
  wire  _T_993; // @[CSR.scala 578:73]
  wire  _T_994; // @[CSR.scala 578:73]
  wire  _T_995; // @[CSR.scala 578:73]
  wire  _T_996; // @[CSR.scala 578:73]
  wire  _T_997; // @[CSR.scala 578:73]
  wire  _T_998; // @[CSR.scala 578:73]
  wire  _T_999; // @[CSR.scala 578:73]
  wire  _T_1087; // @[CSR.scala 578:73]
  wire  _T_1088; // @[CSR.scala 578:73]
  wire  _T_1089; // @[CSR.scala 578:73]
  wire  _T_1090; // @[CSR.scala 578:73]
  wire  _T_1091; // @[CSR.scala 578:73]
  wire  _T_1092; // @[CSR.scala 578:73]
  wire  _T_1093; // @[CSR.scala 578:73]
  wire  _T_1094; // @[CSR.scala 578:73]
  wire  _T_1095; // @[CSR.scala 578:73]
  wire  _T_1096; // @[CSR.scala 578:73]
  wire  _T_1097; // @[CSR.scala 578:73]
  wire  _T_1098; // @[CSR.scala 578:73]
  wire  _T_1099; // @[CSR.scala 578:73]
  wire  _T_1100; // @[CSR.scala 578:73]
  wire  _T_1101; // @[CSR.scala 578:73]
  wire  _T_1102; // @[CSR.scala 578:73]
  wire  _T_1103; // @[CSR.scala 578:73]
  wire  _T_1104; // @[CSR.scala 578:73]
  wire  _T_1105; // @[CSR.scala 578:73]
  wire  _T_1106; // @[CSR.scala 578:73]
  wire  _T_1107; // @[CSR.scala 578:73]
  wire  _T_1109; // @[CSR.scala 578:73]
  wire  _T_1110; // @[CSR.scala 578:73]
  wire  _T_1111; // @[CSR.scala 578:73]
  wire  _T_1112; // @[CSR.scala 578:73]
  wire  _T_1113; // @[CSR.scala 578:73]
  wire  _T_1114; // @[CSR.scala 578:73]
  wire  _T_1115; // @[CSR.scala 578:73]
  wire  _T_1116; // @[CSR.scala 578:73]
  wire  _T_1126; // @[CSR.scala 578:73]
  wire [63:0] _T_1130; // @[CSR.scala 1031:9]
  wire [63:0] _T_1131; // @[CSR.scala 1031:34]
  wire  _T_1134; // @[CSR.scala 1031:59]
  wire [63:0] _T_1135; // @[CSR.scala 1031:49]
  wire [63:0] wdata; // @[CSR.scala 1031:43]
  wire [31:0] _T_1150; // @[Decode.scala 14:65]
  wire  _T_1151; // @[Decode.scala 14:121]
  wire  insn_wfi; // @[CSR.scala 590:159]
  wire [31:0] _T_1161; // @[CSR.scala 593:84]
  wire [31:0] _T_1168; // @[Decode.scala 14:65]
  wire  _T_1169; // @[Decode.scala 14:121]
  wire [31:0] _T_1170; // @[Decode.scala 14:65]
  wire  _T_1171; // @[Decode.scala 14:121]
  wire  _T_1173; // @[Decode.scala 15:30]
  wire [31:0] _T_1174; // @[Decode.scala 14:65]
  wire  _T_1175; // @[Decode.scala 14:121]
  wire [31:0] _T_1177; // @[Decode.scala 14:65]
  wire  _T_1178; // @[Decode.scala 14:121]
  wire  _T_1185; // @[CSR.scala 595:55]
  wire  _T_1188; // @[CSR.scala 595:63]
  wire  _T_1192; // @[CSR.scala 596:70]
  wire  _T_1196; // @[CSR.scala 597:64]
  wire [31:0] _T_1199; // @[CSR.scala 599:67]
  wire  _T_1201; // @[CSR.scala 599:50]
  wire  _T_1202; // @[CSR.scala 600:36]
  wire [31:0] _T_1204; // @[CSR.scala 600:62]
  wire  _T_1206; // @[CSR.scala 600:45]
  wire  _T_1207; // @[CSR.scala 599:83]
  wire  _T_1208; // @[CSR.scala 601:39]
  wire [11:0] _T_1212; // @[Decode.scala 14:65]
  wire  _T_1222; // @[CSR.scala 604:44]
  wire  _T_1223; // @[CSR.scala 594:99]
  wire  _T_1224; // @[CSR.scala 594:99]
  wire  _T_1225; // @[CSR.scala 594:99]
  wire  _T_1226; // @[CSR.scala 594:99]
  wire  _T_1227; // @[CSR.scala 594:99]
  wire  _T_1228; // @[CSR.scala 594:99]
  wire  _T_1229; // @[CSR.scala 594:99]
  wire  _T_1230; // @[CSR.scala 594:99]
  wire  _T_1231; // @[CSR.scala 594:99]
  wire  _T_1232; // @[CSR.scala 594:99]
  wire  _T_1233; // @[CSR.scala 594:99]
  wire  _T_1234; // @[CSR.scala 594:99]
  wire  _T_1235; // @[CSR.scala 594:99]
  wire  _T_1236; // @[CSR.scala 594:99]
  wire  _T_1237; // @[CSR.scala 594:99]
  wire  _T_1238; // @[CSR.scala 594:99]
  wire  _T_1239; // @[CSR.scala 594:99]
  wire  _T_1240; // @[CSR.scala 594:99]
  wire  _T_1241; // @[CSR.scala 594:99]
  wire  _T_1242; // @[CSR.scala 594:99]
  wire  _T_1243; // @[CSR.scala 594:99]
  wire  _T_1244; // @[CSR.scala 594:99]
  wire  _T_1245; // @[CSR.scala 594:99]
  wire  _T_1246; // @[CSR.scala 594:99]
  wire  _T_1247; // @[CSR.scala 594:99]
  wire  _T_1248; // @[CSR.scala 594:99]
  wire  _T_1249; // @[CSR.scala 594:99]
  wire  _T_1250; // @[CSR.scala 594:99]
  wire  _T_1251; // @[CSR.scala 594:99]
  wire  _T_1252; // @[CSR.scala 594:99]
  wire  _T_1253; // @[CSR.scala 594:99]
  wire  _T_1254; // @[CSR.scala 594:99]
  wire  _T_1255; // @[CSR.scala 594:99]
  wire  _T_1256; // @[CSR.scala 594:99]
  wire  _T_1257; // @[CSR.scala 594:99]
  wire  _T_1258; // @[CSR.scala 594:99]
  wire  _T_1259; // @[CSR.scala 594:99]
  wire  _T_1260; // @[CSR.scala 594:99]
  wire  _T_1261; // @[CSR.scala 594:99]
  wire  _T_1262; // @[CSR.scala 594:99]
  wire  _T_1263; // @[CSR.scala 594:99]
  wire  _T_1264; // @[CSR.scala 594:99]
  wire  _T_1265; // @[CSR.scala 594:99]
  wire  _T_1266; // @[CSR.scala 594:99]
  wire  _T_1267; // @[CSR.scala 594:99]
  wire  _T_1268; // @[CSR.scala 594:99]
  wire  _T_1269; // @[CSR.scala 594:99]
  wire  _T_1270; // @[CSR.scala 594:99]
  wire  _T_1271; // @[CSR.scala 594:99]
  wire  _T_1272; // @[CSR.scala 594:99]
  wire  _T_1273; // @[CSR.scala 594:99]
  wire  _T_1274; // @[CSR.scala 594:99]
  wire  _T_1275; // @[CSR.scala 594:99]
  wire  _T_1276; // @[CSR.scala 594:99]
  wire  _T_1277; // @[CSR.scala 594:99]
  wire  _T_1278; // @[CSR.scala 594:99]
  wire  _T_1279; // @[CSR.scala 594:99]
  wire  _T_1280; // @[CSR.scala 594:99]
  wire  _T_1281; // @[CSR.scala 594:99]
  wire  _T_1282; // @[CSR.scala 594:99]
  wire  _T_1283; // @[CSR.scala 594:99]
  wire  _T_1284; // @[CSR.scala 594:99]
  wire  _T_1285; // @[CSR.scala 594:99]
  wire  _T_1286; // @[CSR.scala 594:99]
  wire  _T_1287; // @[CSR.scala 594:99]
  wire  _T_1288; // @[CSR.scala 594:99]
  wire  _T_1289; // @[CSR.scala 594:99]
  wire  _T_1290; // @[CSR.scala 594:99]
  wire  _T_1291; // @[CSR.scala 594:99]
  wire  _T_1292; // @[CSR.scala 594:99]
  wire  _T_1293; // @[CSR.scala 594:99]
  wire  _T_1294; // @[CSR.scala 594:99]
  wire  _T_1295; // @[CSR.scala 594:99]
  wire  _T_1296; // @[CSR.scala 594:99]
  wire  _T_1297; // @[CSR.scala 594:99]
  wire  _T_1298; // @[CSR.scala 594:99]
  wire  _T_1299; // @[CSR.scala 594:99]
  wire  _T_1300; // @[CSR.scala 594:99]
  wire  _T_1301; // @[CSR.scala 594:99]
  wire  _T_1302; // @[CSR.scala 594:99]
  wire  _T_1303; // @[CSR.scala 594:99]
  wire  _T_1304; // @[CSR.scala 594:99]
  wire  _T_1305; // @[CSR.scala 594:99]
  wire  _T_1306; // @[CSR.scala 594:99]
  wire  _T_1307; // @[CSR.scala 594:99]
  wire  _T_1308; // @[CSR.scala 594:99]
  wire  _T_1309; // @[CSR.scala 594:99]
  wire  _T_1310; // @[CSR.scala 594:99]
  wire  _T_1311; // @[CSR.scala 594:99]
  wire  _T_1312; // @[CSR.scala 594:99]
  wire  _T_1313; // @[CSR.scala 594:99]
  wire  _T_1314; // @[CSR.scala 594:99]
  wire  _T_1315; // @[CSR.scala 594:99]
  wire  _T_1316; // @[CSR.scala 594:99]
  wire  _T_1317; // @[CSR.scala 594:99]
  wire  _T_1318; // @[CSR.scala 594:99]
  wire  _T_1319; // @[CSR.scala 594:99]
  wire  _T_1320; // @[CSR.scala 594:99]
  wire  _T_1321; // @[CSR.scala 594:99]
  wire  _T_1322; // @[CSR.scala 594:99]
  wire  _T_1323; // @[CSR.scala 594:99]
  wire  _T_1324; // @[CSR.scala 594:99]
  wire  _T_1325; // @[CSR.scala 594:99]
  wire  _T_1326; // @[CSR.scala 594:99]
  wire  _T_1327; // @[CSR.scala 594:99]
  wire  _T_1328; // @[CSR.scala 594:99]
  wire  _T_1329; // @[CSR.scala 594:99]
  wire  _T_1330; // @[CSR.scala 594:99]
  wire  _T_1331; // @[CSR.scala 594:99]
  wire  _T_1332; // @[CSR.scala 594:99]
  wire  _T_1333; // @[CSR.scala 594:99]
  wire  _T_1334; // @[CSR.scala 594:99]
  wire  _T_1335; // @[CSR.scala 594:99]
  wire  _T_1336; // @[CSR.scala 594:99]
  wire  _T_1337; // @[CSR.scala 594:99]
  wire  _T_1338; // @[CSR.scala 594:99]
  wire  _T_1339; // @[CSR.scala 594:99]
  wire  _T_1340; // @[CSR.scala 594:99]
  wire  _T_1341; // @[CSR.scala 594:99]
  wire  _T_1342; // @[CSR.scala 594:99]
  wire  _T_1343; // @[CSR.scala 594:99]
  wire  _T_1344; // @[CSR.scala 594:99]
  wire  _T_1345; // @[CSR.scala 594:99]
  wire  _T_1346; // @[CSR.scala 594:99]
  wire  _T_1347; // @[CSR.scala 594:99]
  wire  _T_1348; // @[CSR.scala 594:99]
  wire  _T_1349; // @[CSR.scala 594:99]
  wire  _T_1350; // @[CSR.scala 594:99]
  wire  _T_1351; // @[CSR.scala 594:99]
  wire  _T_1352; // @[CSR.scala 594:99]
  wire  _T_1353; // @[CSR.scala 594:99]
  wire  _T_1354; // @[CSR.scala 594:99]
  wire  _T_1355; // @[CSR.scala 594:99]
  wire  _T_1356; // @[CSR.scala 594:99]
  wire  _T_1357; // @[CSR.scala 594:99]
  wire  _T_1358; // @[CSR.scala 594:99]
  wire  _T_1359; // @[CSR.scala 594:99]
  wire  _T_1360; // @[CSR.scala 594:99]
  wire  _T_1361; // @[CSR.scala 594:99]
  wire  _T_1362; // @[CSR.scala 594:99]
  wire  _T_1363; // @[CSR.scala 594:99]
  wire  _T_1364; // @[CSR.scala 594:99]
  wire  _T_1365; // @[CSR.scala 594:99]
  wire  _T_1366; // @[CSR.scala 594:99]
  wire  _T_1367; // @[CSR.scala 594:99]
  wire  _T_1368; // @[CSR.scala 594:99]
  wire  _T_1369; // @[CSR.scala 594:99]
  wire  _T_1370; // @[CSR.scala 594:99]
  wire  _T_1371; // @[CSR.scala 594:99]
  wire  _T_1372; // @[CSR.scala 594:99]
  wire  _T_1373; // @[CSR.scala 594:115]
  wire  _T_1374; // @[CSR.scala 594:115]
  wire  _T_1375; // @[CSR.scala 594:115]
  wire  _T_1376; // @[CSR.scala 594:115]
  wire  _T_1377; // @[CSR.scala 594:115]
  wire  _T_1378; // @[CSR.scala 594:115]
  wire  _T_1379; // @[CSR.scala 594:115]
  wire  _T_1380; // @[CSR.scala 594:115]
  wire  _T_1381; // @[CSR.scala 594:115]
  wire  _T_1382; // @[CSR.scala 594:115]
  wire  _T_1383; // @[CSR.scala 594:115]
  wire  _T_1384; // @[CSR.scala 594:115]
  wire  _T_1385; // @[CSR.scala 594:115]
  wire  _T_1386; // @[CSR.scala 594:115]
  wire  _T_1387; // @[CSR.scala 594:115]
  wire  _T_1388; // @[CSR.scala 594:115]
  wire  _T_1389; // @[CSR.scala 594:115]
  wire  _T_1390; // @[CSR.scala 594:115]
  wire  _T_1391; // @[CSR.scala 594:115]
  wire  _T_1392; // @[CSR.scala 594:115]
  wire  _T_1393; // @[CSR.scala 594:115]
  wire  _T_1394; // @[CSR.scala 594:115]
  wire  _T_1395; // @[CSR.scala 594:115]
  wire  _T_1396; // @[CSR.scala 594:115]
  wire  _T_1397; // @[CSR.scala 594:115]
  wire  _T_1398; // @[CSR.scala 594:115]
  wire  _T_1399; // @[CSR.scala 594:115]
  wire  _T_1400; // @[CSR.scala 594:115]
  wire  _T_1401; // @[CSR.scala 594:115]
  wire  _T_1402; // @[CSR.scala 594:115]
  wire  _T_1403; // @[CSR.scala 594:115]
  wire  _T_1404; // @[CSR.scala 594:115]
  wire  _T_1405; // @[CSR.scala 594:115]
  wire  _T_1406; // @[CSR.scala 594:115]
  wire  _T_1407; // @[CSR.scala 594:115]
  wire  _T_1408; // @[CSR.scala 594:115]
  wire  _T_1409; // @[CSR.scala 594:115]
  wire  _T_1410; // @[CSR.scala 594:115]
  wire  _T_1411; // @[CSR.scala 594:115]
  wire  _T_1412; // @[CSR.scala 594:115]
  wire  _T_1413; // @[CSR.scala 594:115]
  wire  _T_1414; // @[CSR.scala 594:115]
  wire  _T_1415; // @[CSR.scala 594:115]
  wire  _T_1416; // @[CSR.scala 594:115]
  wire  _T_1417; // @[CSR.scala 594:115]
  wire  _T_1418; // @[CSR.scala 594:115]
  wire  _T_1419; // @[CSR.scala 594:115]
  wire  _T_1420; // @[CSR.scala 594:115]
  wire  _T_1421; // @[CSR.scala 594:115]
  wire  _T_1422; // @[CSR.scala 594:115]
  wire  _T_1423; // @[CSR.scala 594:115]
  wire  _T_1424; // @[CSR.scala 594:115]
  wire  _T_1425; // @[CSR.scala 594:115]
  wire  _T_1426; // @[CSR.scala 594:115]
  wire  _T_1427; // @[CSR.scala 594:115]
  wire  _T_1428; // @[CSR.scala 594:115]
  wire  _T_1429; // @[CSR.scala 594:115]
  wire  _T_1430; // @[CSR.scala 594:115]
  wire  _T_1431; // @[CSR.scala 594:115]
  wire  _T_1432; // @[CSR.scala 594:115]
  wire  _T_1433; // @[CSR.scala 594:115]
  wire  _T_1434; // @[CSR.scala 594:115]
  wire  _T_1435; // @[CSR.scala 594:115]
  wire  _T_1436; // @[CSR.scala 594:115]
  wire  _T_1437; // @[CSR.scala 594:115]
  wire  _T_1438; // @[CSR.scala 594:115]
  wire  _T_1439; // @[CSR.scala 594:115]
  wire  _T_1440; // @[CSR.scala 594:115]
  wire  _T_1441; // @[CSR.scala 594:115]
  wire  _T_1442; // @[CSR.scala 594:115]
  wire  _T_1443; // @[CSR.scala 594:115]
  wire  _T_1444; // @[CSR.scala 594:115]
  wire  _T_1445; // @[CSR.scala 594:115]
  wire  _T_1446; // @[CSR.scala 594:115]
  wire  _T_1447; // @[CSR.scala 594:115]
  wire  _T_1448; // @[CSR.scala 594:115]
  wire  _T_1449; // @[CSR.scala 594:115]
  wire  _T_1450; // @[CSR.scala 594:115]
  wire  _T_1451; // @[CSR.scala 594:115]
  wire  _T_1452; // @[CSR.scala 594:115]
  wire  _T_1453; // @[CSR.scala 594:115]
  wire  _T_1454; // @[CSR.scala 594:115]
  wire  _T_1455; // @[CSR.scala 594:115]
  wire  _T_1456; // @[CSR.scala 594:115]
  wire  _T_1457; // @[CSR.scala 594:115]
  wire  _T_1458; // @[CSR.scala 594:115]
  wire  _T_1459; // @[CSR.scala 594:115]
  wire  _T_1460; // @[CSR.scala 594:115]
  wire  _T_1461; // @[CSR.scala 594:115]
  wire  _T_1462; // @[CSR.scala 594:115]
  wire  _T_1463; // @[CSR.scala 594:115]
  wire  _T_1464; // @[CSR.scala 594:115]
  wire  _T_1465; // @[CSR.scala 594:115]
  wire  _T_1466; // @[CSR.scala 594:115]
  wire  _T_1467; // @[CSR.scala 594:115]
  wire  _T_1468; // @[CSR.scala 594:115]
  wire  _T_1469; // @[CSR.scala 594:115]
  wire  _T_1470; // @[CSR.scala 594:115]
  wire  _T_1471; // @[CSR.scala 594:115]
  wire  _T_1472; // @[CSR.scala 594:115]
  wire  _T_1473; // @[CSR.scala 594:115]
  wire  _T_1474; // @[CSR.scala 594:115]
  wire  _T_1475; // @[CSR.scala 594:115]
  wire  _T_1476; // @[CSR.scala 594:115]
  wire  _T_1477; // @[CSR.scala 594:115]
  wire  _T_1478; // @[CSR.scala 594:115]
  wire  _T_1479; // @[CSR.scala 594:115]
  wire  _T_1480; // @[CSR.scala 594:115]
  wire  _T_1481; // @[CSR.scala 594:115]
  wire  _T_1482; // @[CSR.scala 594:115]
  wire  _T_1483; // @[CSR.scala 594:115]
  wire  _T_1484; // @[CSR.scala 594:115]
  wire  _T_1485; // @[CSR.scala 594:115]
  wire  _T_1486; // @[CSR.scala 594:115]
  wire  _T_1487; // @[CSR.scala 594:115]
  wire  _T_1488; // @[CSR.scala 594:115]
  wire  _T_1489; // @[CSR.scala 594:115]
  wire  _T_1490; // @[CSR.scala 594:115]
  wire  _T_1491; // @[CSR.scala 594:115]
  wire  _T_1492; // @[CSR.scala 594:115]
  wire  _T_1493; // @[CSR.scala 594:115]
  wire  _T_1494; // @[CSR.scala 594:115]
  wire  _T_1495; // @[CSR.scala 594:115]
  wire  _T_1496; // @[CSR.scala 594:115]
  wire  _T_1497; // @[CSR.scala 594:115]
  wire  _T_1498; // @[CSR.scala 594:115]
  wire  _T_1499; // @[CSR.scala 594:115]
  wire  _T_1500; // @[CSR.scala 594:115]
  wire  _T_1501; // @[CSR.scala 594:115]
  wire  _T_1502; // @[CSR.scala 594:115]
  wire  _T_1503; // @[CSR.scala 594:115]
  wire  _T_1504; // @[CSR.scala 594:115]
  wire  _T_1505; // @[CSR.scala 594:115]
  wire  _T_1506; // @[CSR.scala 594:115]
  wire  _T_1507; // @[CSR.scala 594:115]
  wire  _T_1508; // @[CSR.scala 594:115]
  wire  _T_1509; // @[CSR.scala 594:115]
  wire  _T_1510; // @[CSR.scala 594:115]
  wire  _T_1511; // @[CSR.scala 594:115]
  wire  _T_1512; // @[CSR.scala 594:115]
  wire  _T_1513; // @[CSR.scala 594:115]
  wire  _T_1514; // @[CSR.scala 594:115]
  wire  _T_1515; // @[CSR.scala 594:115]
  wire  _T_1516; // @[CSR.scala 594:115]
  wire  _T_1517; // @[CSR.scala 594:115]
  wire  _T_1518; // @[CSR.scala 594:115]
  wire  _T_1519; // @[CSR.scala 594:115]
  wire  _T_1520; // @[CSR.scala 594:115]
  wire  _T_1521; // @[CSR.scala 594:115]
  wire  _T_1523; // @[CSR.scala 604:62]
  wire  _T_1526; // @[CSR.scala 606:33]
  wire  _T_1527; // @[CSR.scala 605:32]
  wire  _T_1528; // @[package.scala 158:47]
  wire  _T_1529; // @[package.scala 158:60]
  wire  _T_1530; // @[package.scala 158:55]
  wire  _T_1531; // @[package.scala 158:47]
  wire  _T_1532; // @[package.scala 158:60]
  wire  _T_1533; // @[package.scala 158:55]
  wire  _T_1534; // @[CSR.scala 607:66]
  wire  _T_1536; // @[CSR.scala 607:130]
  wire  _T_1537; // @[CSR.scala 606:54]
  wire  _T_1541; // @[CSR.scala 594:115]
  wire  _T_1542; // @[CSR.scala 594:115]
  wire  _T_1545; // @[CSR.scala 608:49]
  wire  _T_1546; // @[CSR.scala 607:148]
  wire  _T_1547; // @[CSR.scala 609:21]
  wire  _T_1552; // @[CSR.scala 611:40]
  wire  _T_1553; // @[CSR.scala 611:71]
  wire  _T_1554; // @[CSR.scala 611:57]
  wire  _T_1555; // @[CSR.scala 611:102]
  wire  _T_1556; // @[CSR.scala 611:133]
  wire  _T_1557; // @[CSR.scala 611:119]
  wire  _T_1558; // @[CSR.scala 611:88]
  wire  _T_1563; // @[CSR.scala 613:14]
  wire  _T_1564; // @[CSR.scala 612:64]
  wire  _T_1566; // @[CSR.scala 614:14]
  wire  _T_1567; // @[CSR.scala 613:28]
  wire  _T_1569; // @[CSR.scala 615:17]
  wire [11:0] _T_1591; // @[CSR.scala 626:37]
  wire [11:0] debugTVec; // @[CSR.scala 626:22]
  wire [39:0] _T_1601; // @[Cat.scala 30:58]
  wire [39:0] _T_1602; // @[CSR.scala 634:19]
  wire [7:0] _T_1604; // @[CSR.scala 635:59]
  wire [39:0] _T_1606; // @[Cat.scala 30:58]
  wire  _T_1609; // @[CSR.scala 637:28]
  wire  _T_1611; // @[CSR.scala 637:94]
  wire  _T_1612; // @[CSR.scala 637:55]
  wire [39:0] notDebugTVec; // @[CSR.scala 638:8]
  wire [39:0] tvec; // @[CSR.scala 640:17]
  wire  _T_1618; // @[CSR.scala 646:32]
  wire  _T_1620; // @[CSR.scala 646:53]
  wire  _T_1623; // @[CSR.scala 651:53]
  reg [1:0] _T_1626; // @[CSR.scala 651:24]
  reg [31:0] _RAND_123;
  wire [1:0] _T_1628; // @[Bitwise.scala 48:55]
  wire [1:0] _T_1629; // @[Bitwise.scala 48:55]
  wire [2:0] _T_1630; // @[Bitwise.scala 48:55]
  wire  _T_1631; // @[CSR.scala 656:79]
  wire  _T_1633; // @[CSR.scala 656:9]
  wire  _T_1636; // @[CSR.scala 658:18]
  wire  _T_1638; // @[CSR.scala 658:36]
  wire  _GEN_66; // @[CSR.scala 658:51]
  wire  _T_1639; // @[CSR.scala 659:28]
  wire  _T_1640; // @[CSR.scala 659:32]
  wire  _T_1641; // @[CSR.scala 659:55]
  wire  _T_1643; // @[CSR.scala 661:22]
  wire  _GEN_68; // @[CSR.scala 661:36]
  wire  _T_1653; // @[CSR.scala 664:29]
  wire  _T_1655; // @[CSR.scala 664:9]
  wire [39:0] _T_1658; // @[CSR.scala 1052:31]
  wire [39:0] epc; // @[CSR.scala 1052:26]
  wire [1:0] _T_1661; // @[CSR.scala 675:86]
  wire [1:0] _T_1662; // @[CSR.scala 675:56]
  wire  _GEN_70; // @[CSR.scala 672:25]
  wire [39:0] _GEN_71; // @[CSR.scala 672:25]
  wire [39:0] _GEN_75; // @[CSR.scala 679:27]
  wire  _GEN_79; // @[CSR.scala 679:27]
  wire [1:0] _GEN_80; // @[CSR.scala 679:27]
  wire [39:0] _GEN_83; // @[CSR.scala 679:27]
  wire  _GEN_86; // @[CSR.scala 679:27]
  wire [1:0] _GEN_87; // @[CSR.scala 679:27]
  wire  _GEN_88; // @[CSR.scala 679:27]
  wire [39:0] _GEN_90; // @[CSR.scala 671:24]
  wire [39:0] _GEN_94; // @[CSR.scala 671:24]
  wire  _GEN_98; // @[CSR.scala 671:24]
  wire [1:0] _GEN_99; // @[CSR.scala 671:24]
  wire [39:0] _GEN_101; // @[CSR.scala 671:24]
  wire  _GEN_104; // @[CSR.scala 671:24]
  wire [1:0] _GEN_105; // @[CSR.scala 671:24]
  wire  _GEN_106; // @[CSR.scala 671:24]
  wire [39:0] _GEN_108; // @[CSR.scala 670:20]
  wire [39:0] _GEN_112; // @[CSR.scala 670:20]
  wire  _GEN_116; // @[CSR.scala 670:20]
  wire [1:0] _GEN_117; // @[CSR.scala 670:20]
  wire [39:0] _GEN_119; // @[CSR.scala 670:20]
  wire  _GEN_122; // @[CSR.scala 670:20]
  wire [1:0] _GEN_123; // @[CSR.scala 670:20]
  wire  _GEN_124; // @[CSR.scala 670:20]
  wire [39:0] _GEN_127; // @[CSR.scala 725:53]
  wire  _GEN_132; // @[CSR.scala 719:44]
  wire [1:0] _GEN_133; // @[CSR.scala 719:44]
  wire [39:0] _GEN_135; // @[CSR.scala 719:44]
  wire [1:0] _GEN_142; // @[CSR.scala 718:19]
  wire [63:0] _T_1942; // @[Mux.scala 19:72]
  wire [63:0] _T_1943; // @[Mux.scala 19:72]
  wire [63:0] _T_1944; // @[Mux.scala 19:72]
  wire [63:0] _T_1945; // @[Mux.scala 19:72]
  wire [31:0] _T_1946; // @[Mux.scala 19:72]
  wire [15:0] _T_1947; // @[Mux.scala 19:72]
  wire [63:0] _T_1948; // @[Mux.scala 19:72]
  wire [63:0] _T_1949; // @[Mux.scala 19:72]
  wire [63:0] _T_1950; // @[Mux.scala 19:72]
  wire [63:0] _T_1951; // @[Mux.scala 19:72]
  wire [63:0] _T_1952; // @[Mux.scala 19:72]
  wire [1:0] _T_1953; // @[Mux.scala 19:72]
  wire [31:0] _T_1954; // @[Mux.scala 19:72]
  wire [63:0] _T_1955; // @[Mux.scala 19:72]
  wire [63:0] _T_1956; // @[Mux.scala 19:72]
  wire [4:0] _T_1957; // @[Mux.scala 19:72]
  wire [2:0] _T_1958; // @[Mux.scala 19:72]
  wire [7:0] _T_1959; // @[Mux.scala 19:72]
  wire [63:0] _T_1960; // @[Mux.scala 19:72]
  wire [63:0] _T_1961; // @[Mux.scala 19:72]
  wire [31:0] _T_2049; // @[Mux.scala 19:72]
  wire [63:0] _T_2050; // @[Mux.scala 19:72]
  wire [63:0] _T_2051; // @[Mux.scala 19:72]
  wire [26:0] _T_2052; // @[Mux.scala 19:72]
  wire [31:0] _T_2053; // @[Mux.scala 19:72]
  wire [31:0] _T_2054; // @[Mux.scala 19:72]
  wire [31:0] _T_2055; // @[Mux.scala 19:72]
  wire [31:0] _T_2056; // @[Mux.scala 19:72]
  wire [63:0] _T_2057; // @[Mux.scala 19:72]
  wire [63:0] _T_2058; // @[Mux.scala 19:72]
  wire [63:0] _T_2059; // @[Mux.scala 19:72]
  wire [63:0] _T_2060; // @[Mux.scala 19:72]
  wire [63:0] _T_2061; // @[Mux.scala 19:72]
  wire [63:0] _T_2062; // @[Mux.scala 19:72]
  wire [63:0] _T_2063; // @[Mux.scala 19:72]
  wire [63:0] _T_2064; // @[Mux.scala 19:72]
  wire [63:0] _T_2065; // @[Mux.scala 19:72]
  wire [31:0] _T_2066; // @[Mux.scala 19:72]
  wire [63:0] _T_2067; // @[Mux.scala 19:72]
  wire [63:0] _T_2068; // @[Mux.scala 19:72]
  wire [63:0] _T_2069; // @[Mux.scala 19:72]
  wire [29:0] _T_2071; // @[Mux.scala 19:72]
  wire [29:0] _T_2072; // @[Mux.scala 19:72]
  wire [29:0] _T_2073; // @[Mux.scala 19:72]
  wire [29:0] _T_2074; // @[Mux.scala 19:72]
  wire [29:0] _T_2075; // @[Mux.scala 19:72]
  wire [29:0] _T_2076; // @[Mux.scala 19:72]
  wire [29:0] _T_2077; // @[Mux.scala 19:72]
  wire [29:0] _T_2078; // @[Mux.scala 19:72]
  wire [63:0] _T_2088; // @[Mux.scala 19:72]
  wire [63:0] _T_2092; // @[Mux.scala 19:72]
  wire [63:0] _T_2093; // @[Mux.scala 19:72]
  wire [63:0] _T_2094; // @[Mux.scala 19:72]
  wire [63:0] _GEN_743; // @[Mux.scala 19:72]
  wire [63:0] _T_2095; // @[Mux.scala 19:72]
  wire [63:0] _GEN_744; // @[Mux.scala 19:72]
  wire [63:0] _T_2096; // @[Mux.scala 19:72]
  wire [63:0] _T_2097; // @[Mux.scala 19:72]
  wire [63:0] _T_2098; // @[Mux.scala 19:72]
  wire [63:0] _T_2099; // @[Mux.scala 19:72]
  wire [63:0] _T_2100; // @[Mux.scala 19:72]
  wire [63:0] _T_2101; // @[Mux.scala 19:72]
  wire [63:0] _GEN_745; // @[Mux.scala 19:72]
  wire [63:0] _T_2102; // @[Mux.scala 19:72]
  wire [63:0] _GEN_746; // @[Mux.scala 19:72]
  wire [63:0] _T_2103; // @[Mux.scala 19:72]
  wire [63:0] _T_2104; // @[Mux.scala 19:72]
  wire [63:0] _T_2105; // @[Mux.scala 19:72]
  wire [63:0] _GEN_747; // @[Mux.scala 19:72]
  wire [63:0] _T_2106; // @[Mux.scala 19:72]
  wire [63:0] _GEN_748; // @[Mux.scala 19:72]
  wire [63:0] _T_2107; // @[Mux.scala 19:72]
  wire [63:0] _GEN_749; // @[Mux.scala 19:72]
  wire [63:0] _T_2108; // @[Mux.scala 19:72]
  wire [63:0] _T_2109; // @[Mux.scala 19:72]
  wire [63:0] _T_2110; // @[Mux.scala 19:72]
  wire [63:0] _GEN_750; // @[Mux.scala 19:72]
  wire [63:0] _T_2198; // @[Mux.scala 19:72]
  wire [63:0] _T_2199; // @[Mux.scala 19:72]
  wire [63:0] _T_2200; // @[Mux.scala 19:72]
  wire [63:0] _GEN_751; // @[Mux.scala 19:72]
  wire [63:0] _T_2201; // @[Mux.scala 19:72]
  wire [63:0] _GEN_752; // @[Mux.scala 19:72]
  wire [63:0] _T_2202; // @[Mux.scala 19:72]
  wire [63:0] _GEN_753; // @[Mux.scala 19:72]
  wire [63:0] _T_2203; // @[Mux.scala 19:72]
  wire [63:0] _GEN_754; // @[Mux.scala 19:72]
  wire [63:0] _T_2204; // @[Mux.scala 19:72]
  wire [63:0] _GEN_755; // @[Mux.scala 19:72]
  wire [63:0] _T_2205; // @[Mux.scala 19:72]
  wire [63:0] _T_2206; // @[Mux.scala 19:72]
  wire [63:0] _T_2207; // @[Mux.scala 19:72]
  wire [63:0] _T_2208; // @[Mux.scala 19:72]
  wire [63:0] _T_2209; // @[Mux.scala 19:72]
  wire [63:0] _T_2210; // @[Mux.scala 19:72]
  wire [63:0] _T_2211; // @[Mux.scala 19:72]
  wire [63:0] _T_2212; // @[Mux.scala 19:72]
  wire [63:0] _T_2213; // @[Mux.scala 19:72]
  wire [63:0] _T_2214; // @[Mux.scala 19:72]
  wire [63:0] _GEN_756; // @[Mux.scala 19:72]
  wire [63:0] _T_2215; // @[Mux.scala 19:72]
  wire [63:0] _T_2216; // @[Mux.scala 19:72]
  wire [63:0] _T_2217; // @[Mux.scala 19:72]
  wire [63:0] _T_2218; // @[Mux.scala 19:72]
  wire [63:0] _GEN_757; // @[Mux.scala 19:72]
  wire [63:0] _T_2220; // @[Mux.scala 19:72]
  wire [63:0] _GEN_758; // @[Mux.scala 19:72]
  wire [63:0] _T_2221; // @[Mux.scala 19:72]
  wire [63:0] _GEN_759; // @[Mux.scala 19:72]
  wire [63:0] _T_2222; // @[Mux.scala 19:72]
  wire [63:0] _GEN_760; // @[Mux.scala 19:72]
  wire [63:0] _T_2223; // @[Mux.scala 19:72]
  wire [63:0] _GEN_761; // @[Mux.scala 19:72]
  wire [63:0] _T_2224; // @[Mux.scala 19:72]
  wire [63:0] _GEN_762; // @[Mux.scala 19:72]
  wire [63:0] _T_2225; // @[Mux.scala 19:72]
  wire [63:0] _GEN_763; // @[Mux.scala 19:72]
  wire [63:0] _T_2226; // @[Mux.scala 19:72]
  wire [63:0] _GEN_764; // @[Mux.scala 19:72]
  wire [63:0] _T_2227; // @[Mux.scala 19:72]
  wire  _T_2242; // @[package.scala 14:47]
  wire  _T_2243; // @[package.scala 14:47]
  wire  _T_2244; // @[package.scala 14:47]
  wire [4:0] _T_3593; // @[CSR.scala 764:30]
  wire [4:0] _GEN_149; // @[CSR.scala 763:30]
  wire  _T_3597; // @[package.scala 14:62]
  wire  csr_wen; // @[package.scala 14:62]
  wire [8:0] _GEN_175; // @[CSR.scala 796:34]
  wire [19:0] _GEN_176; // @[CSR.scala 796:34]
  wire [9:0] _GEN_177; // @[CSR.scala 796:34]
  wire  _GEN_178; // @[CSR.scala 796:34]
  wire  _GEN_179; // @[CSR.scala 796:34]
  wire  _GEN_184; // @[CSR.scala 792:40]
  wire [8:0] _GEN_185; // @[CSR.scala 792:40]
  wire [19:0] _GEN_186; // @[CSR.scala 792:40]
  wire [9:0] _GEN_187; // @[CSR.scala 792:40]
  wire  _GEN_188; // @[CSR.scala 792:40]
  wire  _GEN_189; // @[CSR.scala 792:40]
  wire  _GEN_214; // @[CSR.scala 796:34]
  wire [8:0] _GEN_215; // @[CSR.scala 796:34]
  wire  _GEN_224; // @[CSR.scala 792:40]
  wire [8:0] _GEN_225; // @[CSR.scala 792:40]
  wire  _GEN_254; // @[CSR.scala 796:34]
  wire [8:0] _GEN_255; // @[CSR.scala 796:34]
  wire  _GEN_264; // @[CSR.scala 792:40]
  wire [8:0] _GEN_265; // @[CSR.scala 792:40]
  wire  _GEN_294; // @[CSR.scala 796:34]
  wire [8:0] _GEN_295; // @[CSR.scala 796:34]
  wire  _GEN_304; // @[CSR.scala 792:40]
  wire [8:0] _GEN_305; // @[CSR.scala 792:40]
  wire [100:0] _T_3676;
  wire  _T_3706; // @[CSR.scala 1035:27]
  wire  _T_3708; // @[CSR.scala 1055:73]
  wire [1:0] _GEN_320; // @[CSR.scala 814:39]
  wire  _T_3716; // @[CSR.scala 841:43]
  wire [3:0] _T_3719; // @[CSR.scala 843:38]
  wire [63:0] _GEN_765; // @[CSR.scala 843:32]
  wire [63:0] _T_3720; // @[CSR.scala 843:32]
  wire [63:0] _T_3722; // @[CSR.scala 843:55]
  wire [63:0] _T_3724; // @[CSR.scala 843:73]
  wire [63:0] _T_3725; // @[CSR.scala 843:62]
  wire [15:0] _T_3740; // @[CSR.scala 851:59]
  wire [15:0] _T_3742; // @[CSR.scala 1031:9]
  wire [63:0] _GEN_766; // @[CSR.scala 1031:34]
  wire [63:0] _T_3743; // @[CSR.scala 1031:34]
  wire [63:0] _T_3749; // @[CSR.scala 1031:43]
  wire [63:0] _T_3777; // @[CSR.scala 858:59]
  wire [63:0] _T_3779; // @[CSR.scala 1052:31]
  wire [63:0] _GEN_333; // @[CSR.scala 859:40]
  wire [63:0] _T_3782; // @[CSR.scala 862:64]
  wire [7:0] _T_3784; // @[CSR.scala 862:75]
  wire [63:0] _GEN_767; // @[CSR.scala 862:70]
  wire [63:0] _T_3785; // @[CSR.scala 862:70]
  wire [63:0] _GEN_335; // @[CSR.scala 862:40]
  wire [63:0] _T_3787; // @[CSR.scala 863:62]
  wire [63:0] _GEN_338; // @[CSR.scala 1049:31]
  wire [63:0] _GEN_340; // @[CSR.scala 1049:31]
  wire [63:0] _GEN_343; // @[CSR.scala 876:40]
  wire [63:0] _GEN_345; // @[CSR.scala 877:40]
  wire [63:0] _GEN_347; // @[CSR.scala 878:40]
  wire [63:0] _GEN_348; // @[CSR.scala 878:40]
  wire  _T_3813; // @[CSR.scala 1035:27]
  wire [63:0] _GEN_354; // @[CSR.scala 889:42]
  wire [1:0] _GEN_358; // @[CSR.scala 893:41]
  wire [63:0] _T_3859; // @[CSR.scala 904:52]
  wire [63:0] _T_3860; // @[CSR.scala 904:77]
  wire [63:0] _T_3861; // @[CSR.scala 904:68]
  wire  _T_3894; // @[CSR.scala 910:30]
  wire  _T_3895; // @[CSR.scala 911:30]
  wire  _T_3898; // @[CSR.scala 912:36]
  wire [63:0] _T_3901; // @[CSR.scala 917:64]
  wire [63:0] _T_3903; // @[CSR.scala 917:80]
  wire [63:0] _GEN_370; // @[CSR.scala 919:42]
  wire [63:0] _GEN_371; // @[CSR.scala 920:42]
  wire [63:0] _T_3913; // @[CSR.scala 921:64]
  wire [63:0] _T_3915; // @[CSR.scala 923:65]
  wire [63:0] _T_3916; // @[CSR.scala 924:65]
  wire [63:0] _T_3917; // @[CSR.scala 925:70]
  wire [63:0] _GEN_376; // @[CSR.scala 925:44]
  wire [63:0] _GEN_377; // @[CSR.scala 928:44]
  wire  _T_3921; // @[CSR.scala 934:31]
  wire  _T_3942; // @[CSR.scala 937:36]
  wire  _T_3943; // @[CSR.scala 940:38]
  wire  _T_3945; // @[CSR.scala 947:57]
  wire  _T_3961; // @[PMP.scala 41:20]
  wire  _T_3962; // @[PMP.scala 43:62]
  wire  _T_3963; // @[PMP.scala 43:44]
  wire  _T_3965; // @[CSR.scala 954:45]
  wire [63:0] _GEN_485; // @[CSR.scala 954:71]
  wire  _T_3967; // @[CSR.scala 947:57]
  wire  _T_3983; // @[PMP.scala 41:20]
  wire  _T_3984; // @[PMP.scala 43:62]
  wire  _T_3985; // @[PMP.scala 43:44]
  wire  _T_3987; // @[CSR.scala 954:45]
  wire [63:0] _GEN_492; // @[CSR.scala 954:71]
  wire  _T_3989; // @[CSR.scala 947:57]
  wire  _T_4005; // @[PMP.scala 41:20]
  wire  _T_4006; // @[PMP.scala 43:62]
  wire  _T_4007; // @[PMP.scala 43:44]
  wire  _T_4009; // @[CSR.scala 954:45]
  wire [63:0] _GEN_499; // @[CSR.scala 954:71]
  wire  _T_4011; // @[CSR.scala 947:57]
  wire  _T_4027; // @[PMP.scala 41:20]
  wire  _T_4028; // @[PMP.scala 43:62]
  wire  _T_4029; // @[PMP.scala 43:44]
  wire  _T_4031; // @[CSR.scala 954:45]
  wire [63:0] _GEN_506; // @[CSR.scala 954:71]
  wire  _T_4033; // @[CSR.scala 947:57]
  wire  _T_4049; // @[PMP.scala 41:20]
  wire  _T_4050; // @[PMP.scala 43:62]
  wire  _T_4051; // @[PMP.scala 43:44]
  wire  _T_4053; // @[CSR.scala 954:45]
  wire [63:0] _GEN_513; // @[CSR.scala 954:71]
  wire  _T_4055; // @[CSR.scala 947:57]
  wire  _T_4071; // @[PMP.scala 41:20]
  wire  _T_4072; // @[PMP.scala 43:62]
  wire  _T_4073; // @[PMP.scala 43:44]
  wire  _T_4075; // @[CSR.scala 954:45]
  wire [63:0] _GEN_520; // @[CSR.scala 954:71]
  wire  _T_4077; // @[CSR.scala 947:57]
  wire  _T_4093; // @[PMP.scala 41:20]
  wire  _T_4094; // @[PMP.scala 43:62]
  wire  _T_4095; // @[PMP.scala 43:44]
  wire  _T_4097; // @[CSR.scala 954:45]
  wire [63:0] _GEN_527; // @[CSR.scala 954:71]
  wire  _T_4099; // @[CSR.scala 947:57]
  wire  _T_4117; // @[PMP.scala 43:44]
  wire  _T_4119; // @[CSR.scala 954:45]
  wire [63:0] _GEN_534; // @[CSR.scala 954:71]
  wire [8:0] _GEN_547; // @[CSR.scala 782:18]
  wire [1:0] _GEN_562; // @[CSR.scala 782:18]
  wire [63:0] _GEN_574; // @[CSR.scala 782:18]
  wire [63:0] _GEN_576; // @[CSR.scala 782:18]
  wire [63:0] _GEN_579; // @[CSR.scala 782:18]
  wire [63:0] _GEN_581; // @[CSR.scala 782:18]
  wire [63:0] _GEN_584; // @[CSR.scala 782:18]
  wire [63:0] _GEN_585; // @[CSR.scala 782:18]
  wire [63:0] _GEN_591; // @[CSR.scala 782:18]
  wire [63:0] _GEN_596; // @[CSR.scala 782:18]
  wire [63:0] _GEN_597; // @[CSR.scala 782:18]
  wire [63:0] _GEN_602; // @[CSR.scala 782:18]
  wire [63:0] _GEN_603; // @[CSR.scala 782:18]
  wire [63:0] _GEN_643; // @[CSR.scala 782:18]
  wire [63:0] _GEN_650; // @[CSR.scala 782:18]
  wire [63:0] _GEN_657; // @[CSR.scala 782:18]
  wire [63:0] _GEN_664; // @[CSR.scala 782:18]
  wire [63:0] _GEN_671; // @[CSR.scala 782:18]
  wire [63:0] _GEN_678; // @[CSR.scala 782:18]
  wire [63:0] _GEN_685; // @[CSR.scala 782:18]
  wire [63:0] _GEN_692; // @[CSR.scala 782:18]
  reg [19:0] CSRFile_state; // @[Register tracking CSRFile state]
  reg [31:0] _RAND_124;
  reg  CSRFile_cov [0:1048575]; // @[Coverage map for CSRFile]
  reg [31:0] _RAND_125;
  wire  CSRFile_cov_read_data; // @[Coverage map for CSRFile]
  wire [19:0] CSRFile_cov_read_addr; // @[Coverage map for CSRFile]
  wire  CSRFile_cov_write_data; // @[Coverage map for CSRFile]
  wire [19:0] CSRFile_cov_write_addr; // @[Coverage map for CSRFile]
  wire  CSRFile_cov_write_mask; // @[Coverage map for CSRFile]
  wire  CSRFile_cov_write_en; // @[Coverage map for CSRFile]
  reg [29:0] CSRFile_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_126;
  wire [15:0] reg_singleStepped_shl;
  wire [19:0] reg_singleStepped_pad;
  wire  reg_debug_shl;
  wire [19:0] reg_debug_pad;
  wire [9:0] reg_pmp_7_cfg_a_shl;
  wire [19:0] reg_pmp_7_cfg_a_pad;
  wire [17:0] reg_dcsr_ebreaku_shl;
  wire [19:0] reg_dcsr_ebreaku_pad;
  wire [13:0] reg_dcsr_ebreaks_shl;
  wire [19:0] reg_dcsr_ebreaks_pad;
  wire [7:0] reg_pmp_6_cfg_l_shl;
  wire [19:0] reg_pmp_6_cfg_l_pad;
  wire [14:0] reg_mstatus_mie_shl;
  wire [19:0] reg_mstatus_mie_pad;
  wire [7:0] reg_pmp_2_cfg_l_shl;
  wire [19:0] reg_pmp_2_cfg_l_pad;
  wire  reg_mstatus_mprv_shl;
  wire [19:0] reg_mstatus_mprv_pad;
  wire [14:0] reg_pmp_0_cfg_l_shl;
  wire [19:0] reg_pmp_0_cfg_l_pad;
  wire [7:0] _T_310_shl;
  wire [19:0] _T_310_pad;
  wire [11:0] reg_pmp_3_cfg_l_shl;
  wire [19:0] reg_pmp_3_cfg_l_pad;
  wire [14:0] reg_mip_stip_shl;
  wire [19:0] reg_mip_stip_pad;
  wire  reg_mip_ssip_shl;
  wire [19:0] reg_mip_ssip_pad;
  wire [19:0] reg_pmp_5_cfg_l_shl;
  wire [19:0] reg_pmp_5_cfg_l_pad;
  wire [6:0] reg_mstatus_spp_shl;
  wire [19:0] reg_mstatus_spp_pad;
  wire [3:0] reg_pmp_4_cfg_l_shl;
  wire [19:0] reg_pmp_4_cfg_l_pad;
  wire [5:0] reg_dcsr_ebreakm_shl;
  wire [19:0] reg_dcsr_ebreakm_pad;
  wire [13:0] reg_mip_seip_shl;
  wire [19:0] reg_mip_seip_pad;
  wire [16:0] reg_pmp_1_cfg_l_shl;
  wire [19:0] reg_pmp_1_cfg_l_pad;
  wire [11:0] reg_bp_0_control_dmode_shl;
  wire [19:0] reg_bp_0_control_dmode_pad;
  wire [7:0] reg_pmp_7_cfg_l_shl;
  wire [19:0] reg_pmp_7_cfg_l_pad;
  wire [3:0] reg_mstatus_prv_shl;
  wire [19:0] reg_mstatus_prv_pad;
  wire [19:0] reg_wfi_shl;
  wire [19:0] reg_wfi_pad;
  wire [3:0] reg_mstatus_sie_shl;
  wire [19:0] reg_mstatus_sie_pad;
  wire [15:0] pcode_regs_0_locked_shl;
  wire [19:0] pcode_regs_0_locked_pad;
  wire [15:0] pcode_regs_1_locked_shl;
  wire [19:0] pcode_regs_1_locked_pad;
  wire [15:0] pcode_regs_2_locked_shl;
  wire [19:0] pcode_regs_2_locked_pad;
  wire [15:0] pcode_regs_3_locked_shl;
  wire [19:0] pcode_regs_3_locked_pad;
  wire [19:0] CSRFile_xor16;
  wire [19:0] CSRFile_xor7;
  wire [19:0] CSRFile_xor17;
  wire [19:0] CSRFile_xor18;
  wire [19:0] CSRFile_xor8;
  wire [19:0] CSRFile_xor3;
  wire [19:0] CSRFile_xor20;
  wire [19:0] CSRFile_xor9;
  wire [19:0] CSRFile_xor21;
  wire [19:0] CSRFile_xor22;
  wire [19:0] CSRFile_xor10;
  wire [19:0] CSRFile_xor4;
  wire [19:0] CSRFile_xor1;
  wire [19:0] CSRFile_xor24;
  wire [19:0] CSRFile_xor11;
  wire [19:0] CSRFile_xor25;
  wire [19:0] CSRFile_xor26;
  wire [19:0] CSRFile_xor12;
  wire [19:0] CSRFile_xor5;
  wire [19:0] CSRFile_xor27;
  wire [19:0] CSRFile_xor28;
  wire [19:0] CSRFile_xor13;
  wire [19:0] CSRFile_xor29;
  wire [19:0] CSRFile_xor30;
  wire [19:0] CSRFile_xor14;
  wire [19:0] CSRFile_xor6;
  wire [19:0] CSRFile_xor2;
  wire [19:0] CSRFile_xor0;
  wire  stopEn0;
  wire  stopEn1;
  wire  CSRFile_or0;
  reg  CSRFile_metaAssert;
  reg [31:0] _RAND_127;
  assign system_insn = io_rw_cmd == 3'h4; // @[CSR.scala 581:31]
  assign _T_1137 = {io_rw_addr, 20'h0}; // @[CSR.scala 590:92]
  assign _T_1144 = _T_1137 & 32'h12400000; // @[Decode.scala 14:65]
  assign _T_1145 = _T_1144 == 32'h10000000; // @[Decode.scala 14:121]
  assign _T_1146 = _T_1137 & 32'h40000000; // @[Decode.scala 14:65]
  assign _T_1147 = _T_1146 == 32'h40000000; // @[Decode.scala 14:121]
  assign _T_1149 = _T_1145 | _T_1147; // @[Decode.scala 15:30]
  assign insn_ret = system_insn & _T_1149; // @[CSR.scala 590:159]
  assign _GEN_125 = io_rw_addr[10] ? reg_dcsr_prv : reg_mstatus_mpp; // @[CSR.scala 725:53]
  assign _GEN_134 = io_rw_addr[9] ? _GEN_125 : {{1'd0}, reg_mstatus_spp}; // @[CSR.scala 719:44]
  assign _T_1138 = _T_1137 & 32'h10100000; // @[Decode.scala 14:65]
  assign _T_1139 = _T_1138 == 32'h0; // @[Decode.scala 14:121]
  assign insn_call = system_insn & _T_1139; // @[CSR.scala 590:159]
  assign _T_1142 = _T_1138 == 32'h100000; // @[Decode.scala 14:121]
  assign insn_break = system_insn & _T_1142; // @[CSR.scala 590:159]
  assign _T_1627 = insn_call | insn_break; // @[CSR.scala 655:29]
  assign exception = _T_1627 | io_exception; // @[CSR.scala 655:43]
  assign _GEN_727 = {{2'd0}, reg_mstatus_prv}; // @[CSR.scala 619:36]
  assign _T_1572 = _GEN_727 + 4'h8; // @[CSR.scala 619:36]
  assign _T_1573 = insn_break ? 64'h3 : io_cause; // @[CSR.scala 620:14]
  assign cause = insn_call ? {{60'd0}, _T_1572} : _T_1573; // @[CSR.scala 619:8]
  assign cause_lsbs = cause[7:0]; // @[CSR.scala 621:25]
  assign _T_1575 = cause_lsbs == 8'he; // @[CSR.scala 622:53]
  assign causeIsDebugInt = cause[63] & _T_1575; // @[CSR.scala 622:39]
  assign _T_1587 = reg_singleStepped | causeIsDebugInt; // @[CSR.scala 625:60]
  assign causeIsDebugTrigger = ~cause[63] & _T_1575; // @[CSR.scala 623:44]
  assign _T_1588 = _T_1587 | causeIsDebugTrigger; // @[CSR.scala 625:79]
  assign _T_1581 = ~cause[63] & insn_break; // @[CSR.scala 624:42]
  assign _T_1584 = {reg_dcsr_ebreakm,1'h0,reg_dcsr_ebreaks,reg_dcsr_ebreaku}; // @[Cat.scala 30:58]
  assign _T_1585 = _T_1584 >> reg_mstatus_prv; // @[CSR.scala 624:134]
  assign causeIsDebugBreak = _T_1581 & _T_1585[0]; // @[CSR.scala 624:56]
  assign _T_1589 = _T_1588 | causeIsDebugBreak; // @[CSR.scala 625:102]
  assign trapToDebug = _T_1589 | reg_debug; // @[CSR.scala 625:123]
  assign _GEN_74 = reg_debug ? reg_mstatus_prv : 2'h3; // @[CSR.scala 672:25]
  assign _T_1592 = reg_mstatus_prv <= 2'h1; // @[CSR.scala 627:51]
  assign _T_1595 = reg_mideleg >> cause_lsbs; // @[CSR.scala 627:93]
  assign _T_1597 = reg_medeleg >> cause_lsbs; // @[CSR.scala 627:118]
  assign _T_1599 = cause[63] ? _T_1595[0] : _T_1597[0]; // @[CSR.scala 627:66]
  assign delegate = _T_1592 & _T_1599; // @[CSR.scala 627:60]
  assign _GEN_82 = delegate ? 2'h1 : 2'h3; // @[CSR.scala 679:27]
  assign _GEN_93 = trapToDebug ? _GEN_74 : _GEN_82; // @[CSR.scala 671:24]
  assign _GEN_111 = exception ? _GEN_93 : reg_mstatus_prv; // @[CSR.scala 670:20]
  assign new_prv = insn_ret ? _GEN_134 : _GEN_111; // @[CSR.scala 718:19]
  assign _T_172 = new_prv == 2'h2; // @[CSR.scala 1035:27]
  assign _GEN_728 = {{5'd0}, io_retire}; // @[Counters.scala 47:33]
  assign _T_287 = _T_286 + _GEN_728; // @[Counters.scala 47:33]
  assign _T_292 = _T_289 + 58'h1; // @[Counters.scala 52:43]
  assign _T_293 = {_T_289,_T_286}; // @[Cat.scala 30:58]
  assign _GEN_729 = {{5'd0}, ~reg_wfi}; // @[Counters.scala 47:33]
  assign _T_297 = _T_296 + _GEN_729; // @[Counters.scala 47:33]
  assign _T_302 = _T_299 + 58'h1; // @[Counters.scala 52:43]
  assign _T_303 = {_T_299,_T_296}; // @[Cat.scala 30:58]
  assign mip_seip = reg_mip_seip | _T_310; // @[CSR.scala 370:57]
  assign _T_318 = {io_interrupts_mtip,1'h0,reg_mip_stip,1'h0,io_interrupts_msip,1'h0,reg_mip_ssip,1'h0}; // @[CSR.scala 372:22]
  assign _T_326 = {4'h0,io_interrupts_meip,1'h0,mip_seip,1'h0,_T_318}; // @[CSR.scala 372:22]
  assign read_mip = _T_326 & 16'haaa; // @[CSR.scala 372:29]
  assign _GEN_730 = {{48'd0}, read_mip}; // @[CSR.scala 375:56]
  assign pending_interrupts = _GEN_730 & reg_mie; // @[CSR.scala 375:56]
  assign d_interrupts = {io_interrupts_debug, 14'h0}; // @[CSR.scala 376:42]
  assign _T_329 = _T_1592 | reg_mstatus_mie; // @[CSR.scala 377:51]
  assign _T_331 = ~pending_interrupts | reg_mideleg; // @[CSR.scala 377:93]
  assign m_interrupts = _T_329 ? ~_T_331 : 64'h0; // @[CSR.scala 377:25]
  assign _T_333 = reg_mstatus_prv < 2'h1; // @[CSR.scala 378:42]
  assign _T_334 = reg_mstatus_prv == 2'h1; // @[CSR.scala 378:70]
  assign _T_335 = _T_334 & reg_mstatus_sie; // @[CSR.scala 378:80]
  assign _T_336 = _T_333 | _T_335; // @[CSR.scala 378:50]
  assign _T_337 = pending_interrupts & reg_mideleg; // @[CSR.scala 378:120]
  assign s_interrupts = _T_336 ? _T_337 : 64'h0; // @[CSR.scala 378:25]
  assign _T_376 = d_interrupts[14] | d_interrupts[13]; // @[CSR.scala 1025:90]
  assign _T_377 = _T_376 | d_interrupts[12]; // @[CSR.scala 1025:90]
  assign _T_378 = _T_377 | d_interrupts[11]; // @[CSR.scala 1025:90]
  assign _T_379 = _T_378 | d_interrupts[3]; // @[CSR.scala 1025:90]
  assign _T_380 = _T_379 | d_interrupts[7]; // @[CSR.scala 1025:90]
  assign _T_381 = _T_380 | d_interrupts[9]; // @[CSR.scala 1025:90]
  assign _T_382 = _T_381 | d_interrupts[1]; // @[CSR.scala 1025:90]
  assign _T_383 = _T_382 | d_interrupts[5]; // @[CSR.scala 1025:90]
  assign _T_384 = _T_383 | d_interrupts[8]; // @[CSR.scala 1025:90]
  assign _T_385 = _T_384 | d_interrupts[0]; // @[CSR.scala 1025:90]
  assign _T_386 = _T_385 | d_interrupts[4]; // @[CSR.scala 1025:90]
  assign _T_387 = _T_386 | m_interrupts[15]; // @[CSR.scala 1025:90]
  assign _T_388 = _T_387 | m_interrupts[14]; // @[CSR.scala 1025:90]
  assign _T_389 = _T_388 | m_interrupts[13]; // @[CSR.scala 1025:90]
  assign _T_390 = _T_389 | m_interrupts[12]; // @[CSR.scala 1025:90]
  assign _T_391 = _T_390 | m_interrupts[11]; // @[CSR.scala 1025:90]
  assign _T_392 = _T_391 | m_interrupts[3]; // @[CSR.scala 1025:90]
  assign _T_393 = _T_392 | m_interrupts[7]; // @[CSR.scala 1025:90]
  assign _T_394 = _T_393 | m_interrupts[9]; // @[CSR.scala 1025:90]
  assign _T_395 = _T_394 | m_interrupts[1]; // @[CSR.scala 1025:90]
  assign _T_396 = _T_395 | m_interrupts[5]; // @[CSR.scala 1025:90]
  assign _T_397 = _T_396 | m_interrupts[8]; // @[CSR.scala 1025:90]
  assign _T_398 = _T_397 | m_interrupts[0]; // @[CSR.scala 1025:90]
  assign _T_399 = _T_398 | m_interrupts[4]; // @[CSR.scala 1025:90]
  assign _T_400 = _T_399 | s_interrupts[15]; // @[CSR.scala 1025:90]
  assign _T_401 = _T_400 | s_interrupts[14]; // @[CSR.scala 1025:90]
  assign _T_402 = _T_401 | s_interrupts[13]; // @[CSR.scala 1025:90]
  assign _T_403 = _T_402 | s_interrupts[12]; // @[CSR.scala 1025:90]
  assign _T_404 = _T_403 | s_interrupts[11]; // @[CSR.scala 1025:90]
  assign _T_405 = _T_404 | s_interrupts[3]; // @[CSR.scala 1025:90]
  assign _T_406 = _T_405 | s_interrupts[7]; // @[CSR.scala 1025:90]
  assign _T_407 = _T_406 | s_interrupts[9]; // @[CSR.scala 1025:90]
  assign _T_408 = _T_407 | s_interrupts[1]; // @[CSR.scala 1025:90]
  assign _T_409 = _T_408 | s_interrupts[5]; // @[CSR.scala 1025:90]
  assign _T_410 = _T_409 | s_interrupts[8]; // @[CSR.scala 1025:90]
  assign _T_411 = _T_410 | s_interrupts[0]; // @[CSR.scala 1025:90]
  assign anyInterrupt = _T_411 | s_interrupts[4]; // @[CSR.scala 1025:90]
  assign _T_450 = s_interrupts[0] ? 3'h0 : 3'h4; // @[Mux.scala 31:69]
  assign _T_451 = s_interrupts[8] ? 4'h8 : {{1'd0}, _T_450}; // @[Mux.scala 31:69]
  assign _T_452 = s_interrupts[5] ? 4'h5 : _T_451; // @[Mux.scala 31:69]
  assign _T_453 = s_interrupts[1] ? 4'h1 : _T_452; // @[Mux.scala 31:69]
  assign _T_454 = s_interrupts[9] ? 4'h9 : _T_453; // @[Mux.scala 31:69]
  assign _T_455 = s_interrupts[7] ? 4'h7 : _T_454; // @[Mux.scala 31:69]
  assign _T_456 = s_interrupts[3] ? 4'h3 : _T_455; // @[Mux.scala 31:69]
  assign _T_457 = s_interrupts[11] ? 4'hb : _T_456; // @[Mux.scala 31:69]
  assign _T_458 = s_interrupts[12] ? 4'hc : _T_457; // @[Mux.scala 31:69]
  assign _T_459 = s_interrupts[13] ? 4'hd : _T_458; // @[Mux.scala 31:69]
  assign _T_460 = s_interrupts[14] ? 4'he : _T_459; // @[Mux.scala 31:69]
  assign _T_461 = s_interrupts[15] ? 4'hf : _T_460; // @[Mux.scala 31:69]
  assign _T_462 = m_interrupts[4] ? 4'h4 : _T_461; // @[Mux.scala 31:69]
  assign _T_463 = m_interrupts[0] ? 4'h0 : _T_462; // @[Mux.scala 31:69]
  assign _T_464 = m_interrupts[8] ? 4'h8 : _T_463; // @[Mux.scala 31:69]
  assign _T_465 = m_interrupts[5] ? 4'h5 : _T_464; // @[Mux.scala 31:69]
  assign _T_466 = m_interrupts[1] ? 4'h1 : _T_465; // @[Mux.scala 31:69]
  assign _T_467 = m_interrupts[9] ? 4'h9 : _T_466; // @[Mux.scala 31:69]
  assign _T_468 = m_interrupts[7] ? 4'h7 : _T_467; // @[Mux.scala 31:69]
  assign _T_469 = m_interrupts[3] ? 4'h3 : _T_468; // @[Mux.scala 31:69]
  assign _T_470 = m_interrupts[11] ? 4'hb : _T_469; // @[Mux.scala 31:69]
  assign _T_471 = m_interrupts[12] ? 4'hc : _T_470; // @[Mux.scala 31:69]
  assign _T_472 = m_interrupts[13] ? 4'hd : _T_471; // @[Mux.scala 31:69]
  assign _T_473 = m_interrupts[14] ? 4'he : _T_472; // @[Mux.scala 31:69]
  assign _T_474 = m_interrupts[15] ? 4'hf : _T_473; // @[Mux.scala 31:69]
  assign _T_475 = d_interrupts[4] ? 4'h4 : _T_474; // @[Mux.scala 31:69]
  assign _T_476 = d_interrupts[0] ? 4'h0 : _T_475; // @[Mux.scala 31:69]
  assign _T_477 = d_interrupts[8] ? 4'h8 : _T_476; // @[Mux.scala 31:69]
  assign _T_478 = d_interrupts[5] ? 4'h5 : _T_477; // @[Mux.scala 31:69]
  assign _T_479 = d_interrupts[1] ? 4'h1 : _T_478; // @[Mux.scala 31:69]
  assign _T_480 = d_interrupts[9] ? 4'h9 : _T_479; // @[Mux.scala 31:69]
  assign _T_481 = d_interrupts[7] ? 4'h7 : _T_480; // @[Mux.scala 31:69]
  assign _T_482 = d_interrupts[3] ? 4'h3 : _T_481; // @[Mux.scala 31:69]
  assign _T_483 = d_interrupts[11] ? 4'hb : _T_482; // @[Mux.scala 31:69]
  assign _T_484 = d_interrupts[12] ? 4'hc : _T_483; // @[Mux.scala 31:69]
  assign _T_485 = d_interrupts[13] ? 4'hd : _T_484; // @[Mux.scala 31:69]
  assign whichInterrupt = d_interrupts[14] ? 4'he : _T_485; // @[Mux.scala 31:69]
  assign _GEN_731 = {{60'd0}, whichInterrupt}; // @[CSR.scala 381:43]
  assign _T_488 = anyInterrupt & ~io_singleStep; // @[CSR.scala 382:33]
  assign _T_489 = _T_488 | reg_singleStepped; // @[CSR.scala 382:51]
  assign _T_495 = {reg_pmp_0_addr,reg_pmp_0_cfg_a[0]}; // @[Cat.scala 30:58]
  assign _T_498 = _T_495 + 31'h1; // @[PMP.scala 52:23]
  assign _T_500 = _T_495 & ~_T_498; // @[PMP.scala 52:14]
  assign _T_501 = {_T_500,2'h3}; // @[Cat.scala 30:58]
  assign _T_505 = {reg_pmp_1_addr,reg_pmp_1_cfg_a[0]}; // @[Cat.scala 30:58]
  assign _T_508 = _T_505 + 31'h1; // @[PMP.scala 52:23]
  assign _T_510 = _T_505 & ~_T_508; // @[PMP.scala 52:14]
  assign _T_511 = {_T_510,2'h3}; // @[Cat.scala 30:58]
  assign _T_515 = {reg_pmp_2_addr,reg_pmp_2_cfg_a[0]}; // @[Cat.scala 30:58]
  assign _T_518 = _T_515 + 31'h1; // @[PMP.scala 52:23]
  assign _T_520 = _T_515 & ~_T_518; // @[PMP.scala 52:14]
  assign _T_521 = {_T_520,2'h3}; // @[Cat.scala 30:58]
  assign _T_525 = {reg_pmp_3_addr,reg_pmp_3_cfg_a[0]}; // @[Cat.scala 30:58]
  assign _T_528 = _T_525 + 31'h1; // @[PMP.scala 52:23]
  assign _T_530 = _T_525 & ~_T_528; // @[PMP.scala 52:14]
  assign _T_531 = {_T_530,2'h3}; // @[Cat.scala 30:58]
  assign _T_535 = {reg_pmp_4_addr,reg_pmp_4_cfg_a[0]}; // @[Cat.scala 30:58]
  assign _T_538 = _T_535 + 31'h1; // @[PMP.scala 52:23]
  assign _T_540 = _T_535 & ~_T_538; // @[PMP.scala 52:14]
  assign _T_541 = {_T_540,2'h3}; // @[Cat.scala 30:58]
  assign _T_545 = {reg_pmp_5_addr,reg_pmp_5_cfg_a[0]}; // @[Cat.scala 30:58]
  assign _T_548 = _T_545 + 31'h1; // @[PMP.scala 52:23]
  assign _T_550 = _T_545 & ~_T_548; // @[PMP.scala 52:14]
  assign _T_551 = {_T_550,2'h3}; // @[Cat.scala 30:58]
  assign _T_555 = {reg_pmp_6_addr,reg_pmp_6_cfg_a[0]}; // @[Cat.scala 30:58]
  assign _T_558 = _T_555 + 31'h1; // @[PMP.scala 52:23]
  assign _T_560 = _T_555 & ~_T_558; // @[PMP.scala 52:14]
  assign _T_561 = {_T_560,2'h3}; // @[Cat.scala 30:58]
  assign _T_565 = {reg_pmp_7_addr,reg_pmp_7_cfg_a[0]}; // @[Cat.scala 30:58]
  assign _T_568 = _T_565 + 31'h1; // @[PMP.scala 52:23]
  assign _T_570 = _T_565 & ~_T_568; // @[PMP.scala 52:14]
  assign _T_571 = {_T_570,2'h3}; // @[Cat.scala 30:58]
  assign _T_578 = {io_status_hpie,io_status_spie,io_status_upie,io_status_mie,io_status_hie,io_status_sie,io_status_uie}; // @[CSR.scala 399:38]
  assign _T_585 = {io_status_mprv,io_status_xs,io_status_fs,io_status_mpp,io_status_hpp,io_status_spp,io_status_mpie,_T_578}; // @[CSR.scala 399:38]
  assign _T_591 = {io_status_sd_rv32,io_status_zero1,io_status_tsr,io_status_tw,io_status_tvm,io_status_mxr,io_status_sum}; // @[CSR.scala 399:38]
  assign _T_600 = {io_status_debug,io_status_isa,io_status_dprv,io_status_prv,io_status_sd,io_status_zero2,io_status_sxl,io_status_uxl,_T_591,_T_585}; // @[CSR.scala 399:38]
  assign read_mstatus = _T_600[63:0]; // @[CSR.scala 399:40]
  assign _T_607 = {reg_bp_0_control_m,1'h0,reg_bp_0_control_s,reg_bp_0_control_u,reg_bp_0_control_x,reg_bp_0_control_w,reg_bp_0_control_r}; // @[CSR.scala 403:48]
  assign _T_615 = {4'h2,reg_bp_0_control_dmode,46'h40000000000,reg_bp_0_control_action,1'h0,2'h0,reg_bp_0_control_tmatch,_T_607}; // @[CSR.scala 403:48]
  assign _T_619 = reg_bp_0_address[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  assign _T_620 = {_T_619,reg_bp_0_address}; // @[Cat.scala 30:58]
  assign _T_623 = reg_misa[2] ? 2'h1 : 2'h3; // @[CSR.scala 1053:36]
  assign _GEN_732 = {{38'd0}, _T_623}; // @[CSR.scala 1053:31]
  assign _T_624 = ~reg_mepc | _GEN_732; // @[CSR.scala 1053:31]
  assign _T_626 = ~_T_624[39]; // @[package.scala 106:38]
  assign _T_628 = _T_626 ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  assign _T_629 = {_T_628,~_T_624}; // @[Cat.scala 30:58]
  assign _T_632 = reg_mbadaddr[39] ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  assign _T_633 = {_T_632,reg_mbadaddr}; // @[Cat.scala 30:58]
  assign _T_639 = {2'h0,1'h0,reg_dcsr_cause,3'h0,reg_dcsr_step,reg_dcsr_prv}; // @[CSR.scala 417:27]
  assign _T_646 = {4'h4,12'h0,reg_dcsr_ebreakm,1'h0,reg_dcsr_ebreaks,reg_dcsr_ebreaku,_T_639}; // @[CSR.scala 417:27]
  assign _T_650 = ~reg_dpc | _GEN_732; // @[CSR.scala 1053:31]
  assign _T_652 = ~_T_650[39]; // @[package.scala 106:38]
  assign _T_654 = _T_652 ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  assign _T_655 = {_T_654,~_T_650}; // @[Cat.scala 30:58]
  assign _T_656 = {reg_frm,reg_fflags}; // @[Cat.scala 30:58]
  assign _T_771 = {30'h0,1'h0,pcode_regs_0_locked}; // @[Cat.scala 30:58]
  assign _T_774 = {30'h0,1'h0,pcode_regs_1_locked}; // @[Cat.scala 30:58]
  assign _T_777 = {30'h0,1'h0,pcode_regs_2_locked}; // @[Cat.scala 30:58]
  assign _T_780 = {30'h0,1'h0,pcode_regs_3_locked}; // @[Cat.scala 30:58]
  assign _T_781 = reg_mie & reg_mideleg; // @[CSR.scala 527:28]
  assign _T_782 = _GEN_730 & reg_mideleg; // @[CSR.scala 528:29]
  assign _T_824 = {1'h0,io_status_spie,2'h0,1'h0,io_status_sie,1'h0}; // @[CSR.scala 541:57]
  assign _T_831 = {1'h0,io_status_xs,io_status_fs,2'h0,2'h0,io_status_spp,1'h0,_T_824}; // @[CSR.scala 541:57]
  assign _T_837 = {io_status_sd_rv32,8'h0,2'h0,1'h0,io_status_mxr,io_status_sum}; // @[CSR.scala 541:57]
  assign _T_846 = {37'h0,io_status_sd,27'h0,2'h0,io_status_uxl,_T_837,_T_831}; // @[CSR.scala 541:57]
  assign _T_850 = reg_sbadaddr[39] ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  assign _T_851 = {_T_850,reg_sbadaddr}; // @[Cat.scala 30:58]
  assign _T_853 = {reg_sptbr_mode,16'h0,reg_sptbr_ppn}; // @[CSR.scala 547:45]
  assign _T_857 = ~reg_sepc | _GEN_732; // @[CSR.scala 1053:31]
  assign _T_859 = ~_T_857[39]; // @[package.scala 106:38]
  assign _T_861 = _T_859 ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  assign _T_862 = {_T_861,~_T_857}; // @[Cat.scala 30:58]
  assign _T_865 = reg_stvec[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  assign _T_866 = {_T_865,reg_stvec}; // @[Cat.scala 30:58]
  assign _T_885 = {reg_pmp_0_cfg_l,2'h0,reg_pmp_0_cfg_a,reg_pmp_0_cfg_x,reg_pmp_0_cfg_w,reg_pmp_0_cfg_r}; // @[package.scala 35:38]
  assign _T_895 = {reg_pmp_2_cfg_l,2'h0,reg_pmp_2_cfg_a,reg_pmp_2_cfg_x,reg_pmp_2_cfg_w,reg_pmp_2_cfg_r}; // @[package.scala 35:38]
  assign _T_905 = {reg_pmp_4_cfg_l,2'h0,reg_pmp_4_cfg_a,reg_pmp_4_cfg_x,reg_pmp_4_cfg_w,reg_pmp_4_cfg_r}; // @[package.scala 35:38]
  assign _T_915 = {reg_pmp_6_cfg_l,2'h0,reg_pmp_6_cfg_a,reg_pmp_6_cfg_x,reg_pmp_6_cfg_w,reg_pmp_6_cfg_r}; // @[package.scala 35:38]
  assign _T_921 = {reg_pmp_1_cfg_l,2'h0,reg_pmp_1_cfg_a,reg_pmp_1_cfg_x,reg_pmp_1_cfg_w,reg_pmp_1_cfg_r,_T_885}; // @[Cat.scala 30:58]
  assign _T_923 = {reg_pmp_3_cfg_l,2'h0,reg_pmp_3_cfg_a,reg_pmp_3_cfg_x,reg_pmp_3_cfg_w,reg_pmp_3_cfg_r,_T_895,_T_921}; // @[Cat.scala 30:58]
  assign _T_924 = {reg_pmp_5_cfg_l,2'h0,reg_pmp_5_cfg_a,reg_pmp_5_cfg_x,reg_pmp_5_cfg_w,reg_pmp_5_cfg_r,_T_905}; // @[Cat.scala 30:58]
  assign _T_927 = {reg_pmp_7_cfg_l,2'h0,reg_pmp_7_cfg_a,reg_pmp_7_cfg_x,reg_pmp_7_cfg_w,reg_pmp_7_cfg_r,_T_915,_T_924,_T_923}; // @[Cat.scala 30:58]
  assign _T_980 = io_rw_addr == 12'h7a1; // @[CSR.scala 578:73]
  assign _T_981 = io_rw_addr == 12'h7a2; // @[CSR.scala 578:73]
  assign _T_982 = io_rw_addr == 12'h301; // @[CSR.scala 578:73]
  assign _T_983 = io_rw_addr == 12'h300; // @[CSR.scala 578:73]
  assign _T_984 = io_rw_addr == 12'h305; // @[CSR.scala 578:73]
  assign _T_985 = io_rw_addr == 12'h344; // @[CSR.scala 578:73]
  assign _T_986 = io_rw_addr == 12'h304; // @[CSR.scala 578:73]
  assign _T_987 = io_rw_addr == 12'h340; // @[CSR.scala 578:73]
  assign _T_988 = io_rw_addr == 12'h341; // @[CSR.scala 578:73]
  assign _T_989 = io_rw_addr == 12'h343; // @[CSR.scala 578:73]
  assign _T_990 = io_rw_addr == 12'h342; // @[CSR.scala 578:73]
  assign _T_991 = io_rw_addr == 12'hf14; // @[CSR.scala 578:73]
  assign _T_992 = io_rw_addr == 12'h7b0; // @[CSR.scala 578:73]
  assign _T_993 = io_rw_addr == 12'h7b1; // @[CSR.scala 578:73]
  assign _T_994 = io_rw_addr == 12'h7b2; // @[CSR.scala 578:73]
  assign _T_995 = io_rw_addr == 12'h1; // @[CSR.scala 578:73]
  assign _T_996 = io_rw_addr == 12'h2; // @[CSR.scala 578:73]
  assign _T_997 = io_rw_addr == 12'h3; // @[CSR.scala 578:73]
  assign _T_998 = io_rw_addr == 12'hb00; // @[CSR.scala 578:73]
  assign _T_999 = io_rw_addr == 12'hb02; // @[CSR.scala 578:73]
  assign _T_1087 = io_rw_addr == 12'h306; // @[CSR.scala 578:73]
  assign _T_1088 = io_rw_addr == 12'hc00; // @[CSR.scala 578:73]
  assign _T_1089 = io_rw_addr == 12'hc02; // @[CSR.scala 578:73]
  assign _T_1090 = io_rw_addr == 12'h182; // @[CSR.scala 578:73]
  assign _T_1091 = io_rw_addr == 12'h190; // @[CSR.scala 578:73]
  assign _T_1092 = io_rw_addr == 12'h191; // @[CSR.scala 578:73]
  assign _T_1093 = io_rw_addr == 12'h192; // @[CSR.scala 578:73]
  assign _T_1094 = io_rw_addr == 12'h193; // @[CSR.scala 578:73]
  assign _T_1095 = io_rw_addr == 12'h100; // @[CSR.scala 578:73]
  assign _T_1096 = io_rw_addr == 12'h144; // @[CSR.scala 578:73]
  assign _T_1097 = io_rw_addr == 12'h104; // @[CSR.scala 578:73]
  assign _T_1098 = io_rw_addr == 12'h140; // @[CSR.scala 578:73]
  assign _T_1099 = io_rw_addr == 12'h142; // @[CSR.scala 578:73]
  assign _T_1100 = io_rw_addr == 12'h143; // @[CSR.scala 578:73]
  assign _T_1101 = io_rw_addr == 12'h180; // @[CSR.scala 578:73]
  assign _T_1102 = io_rw_addr == 12'h141; // @[CSR.scala 578:73]
  assign _T_1103 = io_rw_addr == 12'h105; // @[CSR.scala 578:73]
  assign _T_1104 = io_rw_addr == 12'h106; // @[CSR.scala 578:73]
  assign _T_1105 = io_rw_addr == 12'h303; // @[CSR.scala 578:73]
  assign _T_1106 = io_rw_addr == 12'h302; // @[CSR.scala 578:73]
  assign _T_1107 = io_rw_addr == 12'h3a0; // @[CSR.scala 578:73]
  assign _T_1109 = io_rw_addr == 12'h3b0; // @[CSR.scala 578:73]
  assign _T_1110 = io_rw_addr == 12'h3b1; // @[CSR.scala 578:73]
  assign _T_1111 = io_rw_addr == 12'h3b2; // @[CSR.scala 578:73]
  assign _T_1112 = io_rw_addr == 12'h3b3; // @[CSR.scala 578:73]
  assign _T_1113 = io_rw_addr == 12'h3b4; // @[CSR.scala 578:73]
  assign _T_1114 = io_rw_addr == 12'h3b5; // @[CSR.scala 578:73]
  assign _T_1115 = io_rw_addr == 12'h3b6; // @[CSR.scala 578:73]
  assign _T_1116 = io_rw_addr == 12'h3b7; // @[CSR.scala 578:73]
  assign _T_1126 = io_rw_addr == 12'hf12; // @[CSR.scala 578:73]
  assign _T_1130 = io_rw_cmd[1] ? io_rw_rdata : 64'h0; // @[CSR.scala 1031:9]
  assign _T_1131 = _T_1130 | io_rw_wdata; // @[CSR.scala 1031:34]
  assign _T_1134 = ~io_rw_cmd[1:0] == 2'h0; // @[CSR.scala 1031:59]
  assign _T_1135 = _T_1134 ? io_rw_wdata : 64'h0; // @[CSR.scala 1031:49]
  assign wdata = _T_1131 & ~_T_1135; // @[CSR.scala 1031:43]
  assign _T_1150 = _T_1137 & 32'h12200000; // @[Decode.scala 14:65]
  assign _T_1151 = _T_1150 == 32'h10000000; // @[Decode.scala 14:121]
  assign insn_wfi = system_insn & _T_1151; // @[CSR.scala 590:159]
  assign _T_1161 = {io_decode_0_csr, 20'h0}; // @[CSR.scala 593:84]
  assign _T_1168 = _T_1161 & 32'h12400000; // @[Decode.scala 14:65]
  assign _T_1169 = _T_1168 == 32'h10000000; // @[Decode.scala 14:121]
  assign _T_1170 = _T_1161 & 32'h40000000; // @[Decode.scala 14:65]
  assign _T_1171 = _T_1170 == 32'h40000000; // @[Decode.scala 14:121]
  assign _T_1173 = _T_1169 | _T_1171; // @[Decode.scala 15:30]
  assign _T_1174 = _T_1161 & 32'h12200000; // @[Decode.scala 14:65]
  assign _T_1175 = _T_1174 == 32'h10000000; // @[Decode.scala 14:121]
  assign _T_1177 = _T_1161 & 32'h42000000; // @[Decode.scala 14:65]
  assign _T_1178 = _T_1177 == 32'h2000000; // @[Decode.scala 14:121]
  assign _T_1185 = reg_mstatus_prv > 2'h1; // @[CSR.scala 595:55]
  assign _T_1188 = _T_1185 | ~reg_mstatus_tw; // @[CSR.scala 595:63]
  assign _T_1192 = _T_1185 | ~reg_mstatus_tvm; // @[CSR.scala 596:70]
  assign _T_1196 = _T_1185 | ~reg_mstatus_tsr; // @[CSR.scala 597:64]
  assign _T_1199 = reg_mcounteren >> io_decode_0_csr[4:0]; // @[CSR.scala 599:67]
  assign _T_1201 = _T_1185 | _T_1199[0]; // @[CSR.scala 599:50]
  assign _T_1202 = reg_mstatus_prv >= 2'h1; // @[CSR.scala 600:36]
  assign _T_1204 = reg_scounteren >> io_decode_0_csr[4:0]; // @[CSR.scala 600:62]
  assign _T_1206 = _T_1202 | _T_1204[0]; // @[CSR.scala 600:45]
  assign _T_1207 = _T_1201 & _T_1206; // @[CSR.scala 599:83]
  assign _T_1208 = io_status_fs == 2'h0; // @[CSR.scala 601:39]
  assign _T_1212 = io_decode_0_csr & 12'h900; // @[Decode.scala 14:65]
  assign _T_1222 = reg_mstatus_prv < io_decode_0_csr[9:8]; // @[CSR.scala 604:44]
  assign _T_1223 = io_decode_0_csr == 12'h7a0; // @[CSR.scala 594:99]
  assign _T_1224 = io_decode_0_csr == 12'h7a1; // @[CSR.scala 594:99]
  assign _T_1225 = io_decode_0_csr == 12'h7a2; // @[CSR.scala 594:99]
  assign _T_1226 = io_decode_0_csr == 12'h301; // @[CSR.scala 594:99]
  assign _T_1227 = io_decode_0_csr == 12'h300; // @[CSR.scala 594:99]
  assign _T_1228 = io_decode_0_csr == 12'h305; // @[CSR.scala 594:99]
  assign _T_1229 = io_decode_0_csr == 12'h344; // @[CSR.scala 594:99]
  assign _T_1230 = io_decode_0_csr == 12'h304; // @[CSR.scala 594:99]
  assign _T_1231 = io_decode_0_csr == 12'h340; // @[CSR.scala 594:99]
  assign _T_1232 = io_decode_0_csr == 12'h341; // @[CSR.scala 594:99]
  assign _T_1233 = io_decode_0_csr == 12'h343; // @[CSR.scala 594:99]
  assign _T_1234 = io_decode_0_csr == 12'h342; // @[CSR.scala 594:99]
  assign _T_1235 = io_decode_0_csr == 12'hf14; // @[CSR.scala 594:99]
  assign _T_1236 = io_decode_0_csr == 12'h7b0; // @[CSR.scala 594:99]
  assign _T_1237 = io_decode_0_csr == 12'h7b1; // @[CSR.scala 594:99]
  assign _T_1238 = io_decode_0_csr == 12'h7b2; // @[CSR.scala 594:99]
  assign _T_1239 = io_decode_0_csr == 12'h1; // @[CSR.scala 594:99]
  assign _T_1240 = io_decode_0_csr == 12'h2; // @[CSR.scala 594:99]
  assign _T_1241 = io_decode_0_csr == 12'h3; // @[CSR.scala 594:99]
  assign _T_1242 = io_decode_0_csr == 12'hb00; // @[CSR.scala 594:99]
  assign _T_1243 = io_decode_0_csr == 12'hb02; // @[CSR.scala 594:99]
  assign _T_1244 = io_decode_0_csr == 12'h323; // @[CSR.scala 594:99]
  assign _T_1245 = io_decode_0_csr == 12'hb03; // @[CSR.scala 594:99]
  assign _T_1246 = io_decode_0_csr == 12'hc03; // @[CSR.scala 594:99]
  assign _T_1247 = io_decode_0_csr == 12'h324; // @[CSR.scala 594:99]
  assign _T_1248 = io_decode_0_csr == 12'hb04; // @[CSR.scala 594:99]
  assign _T_1249 = io_decode_0_csr == 12'hc04; // @[CSR.scala 594:99]
  assign _T_1250 = io_decode_0_csr == 12'h325; // @[CSR.scala 594:99]
  assign _T_1251 = io_decode_0_csr == 12'hb05; // @[CSR.scala 594:99]
  assign _T_1252 = io_decode_0_csr == 12'hc05; // @[CSR.scala 594:99]
  assign _T_1253 = io_decode_0_csr == 12'h326; // @[CSR.scala 594:99]
  assign _T_1254 = io_decode_0_csr == 12'hb06; // @[CSR.scala 594:99]
  assign _T_1255 = io_decode_0_csr == 12'hc06; // @[CSR.scala 594:99]
  assign _T_1256 = io_decode_0_csr == 12'h327; // @[CSR.scala 594:99]
  assign _T_1257 = io_decode_0_csr == 12'hb07; // @[CSR.scala 594:99]
  assign _T_1258 = io_decode_0_csr == 12'hc07; // @[CSR.scala 594:99]
  assign _T_1259 = io_decode_0_csr == 12'h328; // @[CSR.scala 594:99]
  assign _T_1260 = io_decode_0_csr == 12'hb08; // @[CSR.scala 594:99]
  assign _T_1261 = io_decode_0_csr == 12'hc08; // @[CSR.scala 594:99]
  assign _T_1262 = io_decode_0_csr == 12'h329; // @[CSR.scala 594:99]
  assign _T_1263 = io_decode_0_csr == 12'hb09; // @[CSR.scala 594:99]
  assign _T_1264 = io_decode_0_csr == 12'hc09; // @[CSR.scala 594:99]
  assign _T_1265 = io_decode_0_csr == 12'h32a; // @[CSR.scala 594:99]
  assign _T_1266 = io_decode_0_csr == 12'hb0a; // @[CSR.scala 594:99]
  assign _T_1267 = io_decode_0_csr == 12'hc0a; // @[CSR.scala 594:99]
  assign _T_1268 = io_decode_0_csr == 12'h32b; // @[CSR.scala 594:99]
  assign _T_1269 = io_decode_0_csr == 12'hb0b; // @[CSR.scala 594:99]
  assign _T_1270 = io_decode_0_csr == 12'hc0b; // @[CSR.scala 594:99]
  assign _T_1271 = io_decode_0_csr == 12'h32c; // @[CSR.scala 594:99]
  assign _T_1272 = io_decode_0_csr == 12'hb0c; // @[CSR.scala 594:99]
  assign _T_1273 = io_decode_0_csr == 12'hc0c; // @[CSR.scala 594:99]
  assign _T_1274 = io_decode_0_csr == 12'h32d; // @[CSR.scala 594:99]
  assign _T_1275 = io_decode_0_csr == 12'hb0d; // @[CSR.scala 594:99]
  assign _T_1276 = io_decode_0_csr == 12'hc0d; // @[CSR.scala 594:99]
  assign _T_1277 = io_decode_0_csr == 12'h32e; // @[CSR.scala 594:99]
  assign _T_1278 = io_decode_0_csr == 12'hb0e; // @[CSR.scala 594:99]
  assign _T_1279 = io_decode_0_csr == 12'hc0e; // @[CSR.scala 594:99]
  assign _T_1280 = io_decode_0_csr == 12'h32f; // @[CSR.scala 594:99]
  assign _T_1281 = io_decode_0_csr == 12'hb0f; // @[CSR.scala 594:99]
  assign _T_1282 = io_decode_0_csr == 12'hc0f; // @[CSR.scala 594:99]
  assign _T_1283 = io_decode_0_csr == 12'h330; // @[CSR.scala 594:99]
  assign _T_1284 = io_decode_0_csr == 12'hb10; // @[CSR.scala 594:99]
  assign _T_1285 = io_decode_0_csr == 12'hc10; // @[CSR.scala 594:99]
  assign _T_1286 = io_decode_0_csr == 12'h331; // @[CSR.scala 594:99]
  assign _T_1287 = io_decode_0_csr == 12'hb11; // @[CSR.scala 594:99]
  assign _T_1288 = io_decode_0_csr == 12'hc11; // @[CSR.scala 594:99]
  assign _T_1289 = io_decode_0_csr == 12'h332; // @[CSR.scala 594:99]
  assign _T_1290 = io_decode_0_csr == 12'hb12; // @[CSR.scala 594:99]
  assign _T_1291 = io_decode_0_csr == 12'hc12; // @[CSR.scala 594:99]
  assign _T_1292 = io_decode_0_csr == 12'h333; // @[CSR.scala 594:99]
  assign _T_1293 = io_decode_0_csr == 12'hb13; // @[CSR.scala 594:99]
  assign _T_1294 = io_decode_0_csr == 12'hc13; // @[CSR.scala 594:99]
  assign _T_1295 = io_decode_0_csr == 12'h334; // @[CSR.scala 594:99]
  assign _T_1296 = io_decode_0_csr == 12'hb14; // @[CSR.scala 594:99]
  assign _T_1297 = io_decode_0_csr == 12'hc14; // @[CSR.scala 594:99]
  assign _T_1298 = io_decode_0_csr == 12'h335; // @[CSR.scala 594:99]
  assign _T_1299 = io_decode_0_csr == 12'hb15; // @[CSR.scala 594:99]
  assign _T_1300 = io_decode_0_csr == 12'hc15; // @[CSR.scala 594:99]
  assign _T_1301 = io_decode_0_csr == 12'h336; // @[CSR.scala 594:99]
  assign _T_1302 = io_decode_0_csr == 12'hb16; // @[CSR.scala 594:99]
  assign _T_1303 = io_decode_0_csr == 12'hc16; // @[CSR.scala 594:99]
  assign _T_1304 = io_decode_0_csr == 12'h337; // @[CSR.scala 594:99]
  assign _T_1305 = io_decode_0_csr == 12'hb17; // @[CSR.scala 594:99]
  assign _T_1306 = io_decode_0_csr == 12'hc17; // @[CSR.scala 594:99]
  assign _T_1307 = io_decode_0_csr == 12'h338; // @[CSR.scala 594:99]
  assign _T_1308 = io_decode_0_csr == 12'hb18; // @[CSR.scala 594:99]
  assign _T_1309 = io_decode_0_csr == 12'hc18; // @[CSR.scala 594:99]
  assign _T_1310 = io_decode_0_csr == 12'h339; // @[CSR.scala 594:99]
  assign _T_1311 = io_decode_0_csr == 12'hb19; // @[CSR.scala 594:99]
  assign _T_1312 = io_decode_0_csr == 12'hc19; // @[CSR.scala 594:99]
  assign _T_1313 = io_decode_0_csr == 12'h33a; // @[CSR.scala 594:99]
  assign _T_1314 = io_decode_0_csr == 12'hb1a; // @[CSR.scala 594:99]
  assign _T_1315 = io_decode_0_csr == 12'hc1a; // @[CSR.scala 594:99]
  assign _T_1316 = io_decode_0_csr == 12'h33b; // @[CSR.scala 594:99]
  assign _T_1317 = io_decode_0_csr == 12'hb1b; // @[CSR.scala 594:99]
  assign _T_1318 = io_decode_0_csr == 12'hc1b; // @[CSR.scala 594:99]
  assign _T_1319 = io_decode_0_csr == 12'h33c; // @[CSR.scala 594:99]
  assign _T_1320 = io_decode_0_csr == 12'hb1c; // @[CSR.scala 594:99]
  assign _T_1321 = io_decode_0_csr == 12'hc1c; // @[CSR.scala 594:99]
  assign _T_1322 = io_decode_0_csr == 12'h33d; // @[CSR.scala 594:99]
  assign _T_1323 = io_decode_0_csr == 12'hb1d; // @[CSR.scala 594:99]
  assign _T_1324 = io_decode_0_csr == 12'hc1d; // @[CSR.scala 594:99]
  assign _T_1325 = io_decode_0_csr == 12'h33e; // @[CSR.scala 594:99]
  assign _T_1326 = io_decode_0_csr == 12'hb1e; // @[CSR.scala 594:99]
  assign _T_1327 = io_decode_0_csr == 12'hc1e; // @[CSR.scala 594:99]
  assign _T_1328 = io_decode_0_csr == 12'h33f; // @[CSR.scala 594:99]
  assign _T_1329 = io_decode_0_csr == 12'hb1f; // @[CSR.scala 594:99]
  assign _T_1330 = io_decode_0_csr == 12'hc1f; // @[CSR.scala 594:99]
  assign _T_1331 = io_decode_0_csr == 12'h306; // @[CSR.scala 594:99]
  assign _T_1332 = io_decode_0_csr == 12'hc00; // @[CSR.scala 594:99]
  assign _T_1333 = io_decode_0_csr == 12'hc02; // @[CSR.scala 594:99]
  assign _T_1334 = io_decode_0_csr == 12'h182; // @[CSR.scala 594:99]
  assign _T_1335 = io_decode_0_csr == 12'h190; // @[CSR.scala 594:99]
  assign _T_1336 = io_decode_0_csr == 12'h191; // @[CSR.scala 594:99]
  assign _T_1337 = io_decode_0_csr == 12'h192; // @[CSR.scala 594:99]
  assign _T_1338 = io_decode_0_csr == 12'h193; // @[CSR.scala 594:99]
  assign _T_1339 = io_decode_0_csr == 12'h100; // @[CSR.scala 594:99]
  assign _T_1340 = io_decode_0_csr == 12'h144; // @[CSR.scala 594:99]
  assign _T_1341 = io_decode_0_csr == 12'h104; // @[CSR.scala 594:99]
  assign _T_1342 = io_decode_0_csr == 12'h140; // @[CSR.scala 594:99]
  assign _T_1343 = io_decode_0_csr == 12'h142; // @[CSR.scala 594:99]
  assign _T_1344 = io_decode_0_csr == 12'h143; // @[CSR.scala 594:99]
  assign _T_1345 = io_decode_0_csr == 12'h180; // @[CSR.scala 594:99]
  assign _T_1346 = io_decode_0_csr == 12'h141; // @[CSR.scala 594:99]
  assign _T_1347 = io_decode_0_csr == 12'h105; // @[CSR.scala 594:99]
  assign _T_1348 = io_decode_0_csr == 12'h106; // @[CSR.scala 594:99]
  assign _T_1349 = io_decode_0_csr == 12'h303; // @[CSR.scala 594:99]
  assign _T_1350 = io_decode_0_csr == 12'h302; // @[CSR.scala 594:99]
  assign _T_1351 = io_decode_0_csr == 12'h3a0; // @[CSR.scala 594:99]
  assign _T_1352 = io_decode_0_csr == 12'h3a2; // @[CSR.scala 594:99]
  assign _T_1353 = io_decode_0_csr == 12'h3b0; // @[CSR.scala 594:99]
  assign _T_1354 = io_decode_0_csr == 12'h3b1; // @[CSR.scala 594:99]
  assign _T_1355 = io_decode_0_csr == 12'h3b2; // @[CSR.scala 594:99]
  assign _T_1356 = io_decode_0_csr == 12'h3b3; // @[CSR.scala 594:99]
  assign _T_1357 = io_decode_0_csr == 12'h3b4; // @[CSR.scala 594:99]
  assign _T_1358 = io_decode_0_csr == 12'h3b5; // @[CSR.scala 594:99]
  assign _T_1359 = io_decode_0_csr == 12'h3b6; // @[CSR.scala 594:99]
  assign _T_1360 = io_decode_0_csr == 12'h3b7; // @[CSR.scala 594:99]
  assign _T_1361 = io_decode_0_csr == 12'h3b8; // @[CSR.scala 594:99]
  assign _T_1362 = io_decode_0_csr == 12'h3b9; // @[CSR.scala 594:99]
  assign _T_1363 = io_decode_0_csr == 12'h3ba; // @[CSR.scala 594:99]
  assign _T_1364 = io_decode_0_csr == 12'h3bb; // @[CSR.scala 594:99]
  assign _T_1365 = io_decode_0_csr == 12'h3bc; // @[CSR.scala 594:99]
  assign _T_1366 = io_decode_0_csr == 12'h3bd; // @[CSR.scala 594:99]
  assign _T_1367 = io_decode_0_csr == 12'h3be; // @[CSR.scala 594:99]
  assign _T_1368 = io_decode_0_csr == 12'h3bf; // @[CSR.scala 594:99]
  assign _T_1369 = io_decode_0_csr == 12'h7c1; // @[CSR.scala 594:99]
  assign _T_1370 = io_decode_0_csr == 12'hf12; // @[CSR.scala 594:99]
  assign _T_1371 = io_decode_0_csr == 12'hf11; // @[CSR.scala 594:99]
  assign _T_1372 = io_decode_0_csr == 12'hf13; // @[CSR.scala 594:99]
  assign _T_1373 = _T_1223 | _T_1224; // @[CSR.scala 594:115]
  assign _T_1374 = _T_1373 | _T_1225; // @[CSR.scala 594:115]
  assign _T_1375 = _T_1374 | _T_1226; // @[CSR.scala 594:115]
  assign _T_1376 = _T_1375 | _T_1227; // @[CSR.scala 594:115]
  assign _T_1377 = _T_1376 | _T_1228; // @[CSR.scala 594:115]
  assign _T_1378 = _T_1377 | _T_1229; // @[CSR.scala 594:115]
  assign _T_1379 = _T_1378 | _T_1230; // @[CSR.scala 594:115]
  assign _T_1380 = _T_1379 | _T_1231; // @[CSR.scala 594:115]
  assign _T_1381 = _T_1380 | _T_1232; // @[CSR.scala 594:115]
  assign _T_1382 = _T_1381 | _T_1233; // @[CSR.scala 594:115]
  assign _T_1383 = _T_1382 | _T_1234; // @[CSR.scala 594:115]
  assign _T_1384 = _T_1383 | _T_1235; // @[CSR.scala 594:115]
  assign _T_1385 = _T_1384 | _T_1236; // @[CSR.scala 594:115]
  assign _T_1386 = _T_1385 | _T_1237; // @[CSR.scala 594:115]
  assign _T_1387 = _T_1386 | _T_1238; // @[CSR.scala 594:115]
  assign _T_1388 = _T_1387 | _T_1239; // @[CSR.scala 594:115]
  assign _T_1389 = _T_1388 | _T_1240; // @[CSR.scala 594:115]
  assign _T_1390 = _T_1389 | _T_1241; // @[CSR.scala 594:115]
  assign _T_1391 = _T_1390 | _T_1242; // @[CSR.scala 594:115]
  assign _T_1392 = _T_1391 | _T_1243; // @[CSR.scala 594:115]
  assign _T_1393 = _T_1392 | _T_1244; // @[CSR.scala 594:115]
  assign _T_1394 = _T_1393 | _T_1245; // @[CSR.scala 594:115]
  assign _T_1395 = _T_1394 | _T_1246; // @[CSR.scala 594:115]
  assign _T_1396 = _T_1395 | _T_1247; // @[CSR.scala 594:115]
  assign _T_1397 = _T_1396 | _T_1248; // @[CSR.scala 594:115]
  assign _T_1398 = _T_1397 | _T_1249; // @[CSR.scala 594:115]
  assign _T_1399 = _T_1398 | _T_1250; // @[CSR.scala 594:115]
  assign _T_1400 = _T_1399 | _T_1251; // @[CSR.scala 594:115]
  assign _T_1401 = _T_1400 | _T_1252; // @[CSR.scala 594:115]
  assign _T_1402 = _T_1401 | _T_1253; // @[CSR.scala 594:115]
  assign _T_1403 = _T_1402 | _T_1254; // @[CSR.scala 594:115]
  assign _T_1404 = _T_1403 | _T_1255; // @[CSR.scala 594:115]
  assign _T_1405 = _T_1404 | _T_1256; // @[CSR.scala 594:115]
  assign _T_1406 = _T_1405 | _T_1257; // @[CSR.scala 594:115]
  assign _T_1407 = _T_1406 | _T_1258; // @[CSR.scala 594:115]
  assign _T_1408 = _T_1407 | _T_1259; // @[CSR.scala 594:115]
  assign _T_1409 = _T_1408 | _T_1260; // @[CSR.scala 594:115]
  assign _T_1410 = _T_1409 | _T_1261; // @[CSR.scala 594:115]
  assign _T_1411 = _T_1410 | _T_1262; // @[CSR.scala 594:115]
  assign _T_1412 = _T_1411 | _T_1263; // @[CSR.scala 594:115]
  assign _T_1413 = _T_1412 | _T_1264; // @[CSR.scala 594:115]
  assign _T_1414 = _T_1413 | _T_1265; // @[CSR.scala 594:115]
  assign _T_1415 = _T_1414 | _T_1266; // @[CSR.scala 594:115]
  assign _T_1416 = _T_1415 | _T_1267; // @[CSR.scala 594:115]
  assign _T_1417 = _T_1416 | _T_1268; // @[CSR.scala 594:115]
  assign _T_1418 = _T_1417 | _T_1269; // @[CSR.scala 594:115]
  assign _T_1419 = _T_1418 | _T_1270; // @[CSR.scala 594:115]
  assign _T_1420 = _T_1419 | _T_1271; // @[CSR.scala 594:115]
  assign _T_1421 = _T_1420 | _T_1272; // @[CSR.scala 594:115]
  assign _T_1422 = _T_1421 | _T_1273; // @[CSR.scala 594:115]
  assign _T_1423 = _T_1422 | _T_1274; // @[CSR.scala 594:115]
  assign _T_1424 = _T_1423 | _T_1275; // @[CSR.scala 594:115]
  assign _T_1425 = _T_1424 | _T_1276; // @[CSR.scala 594:115]
  assign _T_1426 = _T_1425 | _T_1277; // @[CSR.scala 594:115]
  assign _T_1427 = _T_1426 | _T_1278; // @[CSR.scala 594:115]
  assign _T_1428 = _T_1427 | _T_1279; // @[CSR.scala 594:115]
  assign _T_1429 = _T_1428 | _T_1280; // @[CSR.scala 594:115]
  assign _T_1430 = _T_1429 | _T_1281; // @[CSR.scala 594:115]
  assign _T_1431 = _T_1430 | _T_1282; // @[CSR.scala 594:115]
  assign _T_1432 = _T_1431 | _T_1283; // @[CSR.scala 594:115]
  assign _T_1433 = _T_1432 | _T_1284; // @[CSR.scala 594:115]
  assign _T_1434 = _T_1433 | _T_1285; // @[CSR.scala 594:115]
  assign _T_1435 = _T_1434 | _T_1286; // @[CSR.scala 594:115]
  assign _T_1436 = _T_1435 | _T_1287; // @[CSR.scala 594:115]
  assign _T_1437 = _T_1436 | _T_1288; // @[CSR.scala 594:115]
  assign _T_1438 = _T_1437 | _T_1289; // @[CSR.scala 594:115]
  assign _T_1439 = _T_1438 | _T_1290; // @[CSR.scala 594:115]
  assign _T_1440 = _T_1439 | _T_1291; // @[CSR.scala 594:115]
  assign _T_1441 = _T_1440 | _T_1292; // @[CSR.scala 594:115]
  assign _T_1442 = _T_1441 | _T_1293; // @[CSR.scala 594:115]
  assign _T_1443 = _T_1442 | _T_1294; // @[CSR.scala 594:115]
  assign _T_1444 = _T_1443 | _T_1295; // @[CSR.scala 594:115]
  assign _T_1445 = _T_1444 | _T_1296; // @[CSR.scala 594:115]
  assign _T_1446 = _T_1445 | _T_1297; // @[CSR.scala 594:115]
  assign _T_1447 = _T_1446 | _T_1298; // @[CSR.scala 594:115]
  assign _T_1448 = _T_1447 | _T_1299; // @[CSR.scala 594:115]
  assign _T_1449 = _T_1448 | _T_1300; // @[CSR.scala 594:115]
  assign _T_1450 = _T_1449 | _T_1301; // @[CSR.scala 594:115]
  assign _T_1451 = _T_1450 | _T_1302; // @[CSR.scala 594:115]
  assign _T_1452 = _T_1451 | _T_1303; // @[CSR.scala 594:115]
  assign _T_1453 = _T_1452 | _T_1304; // @[CSR.scala 594:115]
  assign _T_1454 = _T_1453 | _T_1305; // @[CSR.scala 594:115]
  assign _T_1455 = _T_1454 | _T_1306; // @[CSR.scala 594:115]
  assign _T_1456 = _T_1455 | _T_1307; // @[CSR.scala 594:115]
  assign _T_1457 = _T_1456 | _T_1308; // @[CSR.scala 594:115]
  assign _T_1458 = _T_1457 | _T_1309; // @[CSR.scala 594:115]
  assign _T_1459 = _T_1458 | _T_1310; // @[CSR.scala 594:115]
  assign _T_1460 = _T_1459 | _T_1311; // @[CSR.scala 594:115]
  assign _T_1461 = _T_1460 | _T_1312; // @[CSR.scala 594:115]
  assign _T_1462 = _T_1461 | _T_1313; // @[CSR.scala 594:115]
  assign _T_1463 = _T_1462 | _T_1314; // @[CSR.scala 594:115]
  assign _T_1464 = _T_1463 | _T_1315; // @[CSR.scala 594:115]
  assign _T_1465 = _T_1464 | _T_1316; // @[CSR.scala 594:115]
  assign _T_1466 = _T_1465 | _T_1317; // @[CSR.scala 594:115]
  assign _T_1467 = _T_1466 | _T_1318; // @[CSR.scala 594:115]
  assign _T_1468 = _T_1467 | _T_1319; // @[CSR.scala 594:115]
  assign _T_1469 = _T_1468 | _T_1320; // @[CSR.scala 594:115]
  assign _T_1470 = _T_1469 | _T_1321; // @[CSR.scala 594:115]
  assign _T_1471 = _T_1470 | _T_1322; // @[CSR.scala 594:115]
  assign _T_1472 = _T_1471 | _T_1323; // @[CSR.scala 594:115]
  assign _T_1473 = _T_1472 | _T_1324; // @[CSR.scala 594:115]
  assign _T_1474 = _T_1473 | _T_1325; // @[CSR.scala 594:115]
  assign _T_1475 = _T_1474 | _T_1326; // @[CSR.scala 594:115]
  assign _T_1476 = _T_1475 | _T_1327; // @[CSR.scala 594:115]
  assign _T_1477 = _T_1476 | _T_1328; // @[CSR.scala 594:115]
  assign _T_1478 = _T_1477 | _T_1329; // @[CSR.scala 594:115]
  assign _T_1479 = _T_1478 | _T_1330; // @[CSR.scala 594:115]
  assign _T_1480 = _T_1479 | _T_1331; // @[CSR.scala 594:115]
  assign _T_1481 = _T_1480 | _T_1332; // @[CSR.scala 594:115]
  assign _T_1482 = _T_1481 | _T_1333; // @[CSR.scala 594:115]
  assign _T_1483 = _T_1482 | _T_1334; // @[CSR.scala 594:115]
  assign _T_1484 = _T_1483 | _T_1335; // @[CSR.scala 594:115]
  assign _T_1485 = _T_1484 | _T_1336; // @[CSR.scala 594:115]
  assign _T_1486 = _T_1485 | _T_1337; // @[CSR.scala 594:115]
  assign _T_1487 = _T_1486 | _T_1338; // @[CSR.scala 594:115]
  assign _T_1488 = _T_1487 | _T_1339; // @[CSR.scala 594:115]
  assign _T_1489 = _T_1488 | _T_1340; // @[CSR.scala 594:115]
  assign _T_1490 = _T_1489 | _T_1341; // @[CSR.scala 594:115]
  assign _T_1491 = _T_1490 | _T_1342; // @[CSR.scala 594:115]
  assign _T_1492 = _T_1491 | _T_1343; // @[CSR.scala 594:115]
  assign _T_1493 = _T_1492 | _T_1344; // @[CSR.scala 594:115]
  assign _T_1494 = _T_1493 | _T_1345; // @[CSR.scala 594:115]
  assign _T_1495 = _T_1494 | _T_1346; // @[CSR.scala 594:115]
  assign _T_1496 = _T_1495 | _T_1347; // @[CSR.scala 594:115]
  assign _T_1497 = _T_1496 | _T_1348; // @[CSR.scala 594:115]
  assign _T_1498 = _T_1497 | _T_1349; // @[CSR.scala 594:115]
  assign _T_1499 = _T_1498 | _T_1350; // @[CSR.scala 594:115]
  assign _T_1500 = _T_1499 | _T_1351; // @[CSR.scala 594:115]
  assign _T_1501 = _T_1500 | _T_1352; // @[CSR.scala 594:115]
  assign _T_1502 = _T_1501 | _T_1353; // @[CSR.scala 594:115]
  assign _T_1503 = _T_1502 | _T_1354; // @[CSR.scala 594:115]
  assign _T_1504 = _T_1503 | _T_1355; // @[CSR.scala 594:115]
  assign _T_1505 = _T_1504 | _T_1356; // @[CSR.scala 594:115]
  assign _T_1506 = _T_1505 | _T_1357; // @[CSR.scala 594:115]
  assign _T_1507 = _T_1506 | _T_1358; // @[CSR.scala 594:115]
  assign _T_1508 = _T_1507 | _T_1359; // @[CSR.scala 594:115]
  assign _T_1509 = _T_1508 | _T_1360; // @[CSR.scala 594:115]
  assign _T_1510 = _T_1509 | _T_1361; // @[CSR.scala 594:115]
  assign _T_1511 = _T_1510 | _T_1362; // @[CSR.scala 594:115]
  assign _T_1512 = _T_1511 | _T_1363; // @[CSR.scala 594:115]
  assign _T_1513 = _T_1512 | _T_1364; // @[CSR.scala 594:115]
  assign _T_1514 = _T_1513 | _T_1365; // @[CSR.scala 594:115]
  assign _T_1515 = _T_1514 | _T_1366; // @[CSR.scala 594:115]
  assign _T_1516 = _T_1515 | _T_1367; // @[CSR.scala 594:115]
  assign _T_1517 = _T_1516 | _T_1368; // @[CSR.scala 594:115]
  assign _T_1518 = _T_1517 | _T_1369; // @[CSR.scala 594:115]
  assign _T_1519 = _T_1518 | _T_1370; // @[CSR.scala 594:115]
  assign _T_1520 = _T_1519 | _T_1371; // @[CSR.scala 594:115]
  assign _T_1521 = _T_1520 | _T_1372; // @[CSR.scala 594:115]
  assign _T_1523 = _T_1222 | ~_T_1521; // @[CSR.scala 604:62]
  assign _T_1526 = _T_1345 & ~_T_1192; // @[CSR.scala 606:33]
  assign _T_1527 = _T_1523 | _T_1526; // @[CSR.scala 605:32]
  assign _T_1528 = io_decode_0_csr >= 12'hc00; // @[package.scala 158:47]
  assign _T_1529 = io_decode_0_csr < 12'hc20; // @[package.scala 158:60]
  assign _T_1530 = _T_1528 & _T_1529; // @[package.scala 158:55]
  assign _T_1531 = io_decode_0_csr >= 12'hc80; // @[package.scala 158:47]
  assign _T_1532 = io_decode_0_csr < 12'hca0; // @[package.scala 158:60]
  assign _T_1533 = _T_1531 & _T_1532; // @[package.scala 158:55]
  assign _T_1534 = _T_1530 | _T_1533; // @[CSR.scala 607:66]
  assign _T_1536 = _T_1534 & ~_T_1207; // @[CSR.scala 607:130]
  assign _T_1537 = _T_1527 | _T_1536; // @[CSR.scala 606:54]
  assign _T_1541 = _T_1236 | _T_1237; // @[CSR.scala 594:115]
  assign _T_1542 = _T_1541 | _T_1238; // @[CSR.scala 594:115]
  assign _T_1545 = _T_1542 & ~reg_debug; // @[CSR.scala 608:49]
  assign _T_1546 = _T_1537 | _T_1545; // @[CSR.scala 607:148]
  assign _T_1547 = io_decode_0_fp_csr & io_decode_0_fp_illegal; // @[CSR.scala 609:21]
  assign _T_1552 = io_decode_0_csr >= 12'h340; // @[CSR.scala 611:40]
  assign _T_1553 = io_decode_0_csr <= 12'h343; // @[CSR.scala 611:71]
  assign _T_1554 = _T_1552 & _T_1553; // @[CSR.scala 611:57]
  assign _T_1555 = io_decode_0_csr >= 12'h140; // @[CSR.scala 611:102]
  assign _T_1556 = io_decode_0_csr <= 12'h143; // @[CSR.scala 611:133]
  assign _T_1557 = _T_1555 & _T_1556; // @[CSR.scala 611:119]
  assign _T_1558 = _T_1554 | _T_1557; // @[CSR.scala 611:88]
  assign _T_1563 = _T_1175 & ~_T_1188; // @[CSR.scala 613:14]
  assign _T_1564 = _T_1222 | _T_1563; // @[CSR.scala 612:64]
  assign _T_1566 = _T_1173 & ~_T_1196; // @[CSR.scala 614:14]
  assign _T_1567 = _T_1564 | _T_1566; // @[CSR.scala 613:28]
  assign _T_1569 = _T_1178 & ~_T_1192; // @[CSR.scala 615:17]
  assign _T_1591 = insn_break ? 12'h800 : 12'h808; // @[CSR.scala 626:37]
  assign debugTVec = reg_debug ? _T_1591 : 12'h800; // @[CSR.scala 626:22]
  assign _T_1601 = {reg_stvec[38],reg_stvec}; // @[Cat.scala 30:58]
  assign _T_1602 = delegate ? _T_1601 : {{8'd0}, reg_mtvec}; // @[CSR.scala 634:19]
  assign _T_1604 = {cause[5:0], 2'h0}; // @[CSR.scala 635:59]
  assign _T_1606 = {_T_1602[39:8],_T_1604}; // @[Cat.scala 30:58]
  assign _T_1609 = _T_1602[0] & cause[63]; // @[CSR.scala 637:28]
  assign _T_1611 = cause_lsbs[7:6] == 2'h0; // @[CSR.scala 637:94]
  assign _T_1612 = _T_1609 & _T_1611; // @[CSR.scala 637:55]
  assign notDebugTVec = _T_1612 ? _T_1606 : _T_1602; // @[CSR.scala 638:8]
  assign tvec = trapToDebug ? {{28'd0}, debugTVec} : notDebugTVec; // @[CSR.scala 640:17]
  assign _T_1618 = ~io_status_fs == 2'h0; // @[CSR.scala 646:32]
  assign _T_1620 = ~io_status_xs == 2'h0; // @[CSR.scala 646:53]
  assign _T_1623 = reg_mstatus_mprv & ~reg_debug; // @[CSR.scala 651:53]
  assign _T_1628 = insn_ret + insn_call; // @[Bitwise.scala 48:55]
  assign _T_1629 = insn_break + io_exception; // @[Bitwise.scala 48:55]
  assign _T_1630 = _T_1628 + _T_1629; // @[Bitwise.scala 48:55]
  assign _T_1631 = _T_1630 <= 3'h1; // @[CSR.scala 656:79]
  assign _T_1633 = _T_1631 | reset; // @[CSR.scala 656:9]
  assign _T_1636 = insn_wfi & ~io_singleStep; // @[CSR.scala 658:18]
  assign _T_1638 = _T_1636 & ~reg_debug; // @[CSR.scala 658:36]
  assign _GEN_66 = _T_1638 | reg_wfi; // @[CSR.scala 658:51]
  assign _T_1639 = pending_interrupts != 64'h0; // @[CSR.scala 659:28]
  assign _T_1640 = _T_1639 | io_interrupts_debug; // @[CSR.scala 659:32]
  assign _T_1641 = _T_1640 | exception; // @[CSR.scala 659:55]
  assign _T_1643 = io_retire | exception; // @[CSR.scala 661:22]
  assign _GEN_68 = _T_1643 | reg_singleStepped; // @[CSR.scala 661:36]
  assign _T_1653 = ~reg_singleStepped | ~io_retire; // @[CSR.scala 664:29]
  assign _T_1655 = _T_1653 | reset; // @[CSR.scala 664:9]
  assign _T_1658 = ~io_pc | 40'h1; // @[CSR.scala 1052:31]
  assign epc = ~_T_1658; // @[CSR.scala 1052:26]
  assign _T_1661 = causeIsDebugTrigger ? 2'h2 : 2'h1; // @[CSR.scala 675:86]
  assign _T_1662 = causeIsDebugInt ? 2'h3 : _T_1661; // @[CSR.scala 675:56]
  assign _GEN_70 = ~reg_debug | reg_debug; // @[CSR.scala 672:25]
  assign _GEN_71 = reg_debug ? reg_dpc : epc; // @[CSR.scala 672:25]
  assign _GEN_75 = delegate ? epc : reg_sepc; // @[CSR.scala 679:27]
  assign _GEN_79 = delegate ? reg_mstatus_sie : reg_mstatus_spie; // @[CSR.scala 679:27]
  assign _GEN_80 = delegate ? reg_mstatus_prv : {{1'd0}, reg_mstatus_spp}; // @[CSR.scala 679:27]
  assign _GEN_83 = delegate ? reg_mepc : epc; // @[CSR.scala 679:27]
  assign _GEN_86 = delegate ? reg_mstatus_mpie : reg_mstatus_mie; // @[CSR.scala 679:27]
  assign _GEN_87 = delegate ? reg_mstatus_mpp : reg_mstatus_prv; // @[CSR.scala 679:27]
  assign _GEN_88 = delegate & reg_mstatus_mie; // @[CSR.scala 679:27]
  assign _GEN_90 = trapToDebug ? _GEN_71 : reg_dpc; // @[CSR.scala 671:24]
  assign _GEN_94 = trapToDebug ? reg_sepc : _GEN_75; // @[CSR.scala 671:24]
  assign _GEN_98 = trapToDebug ? reg_mstatus_spie : _GEN_79; // @[CSR.scala 671:24]
  assign _GEN_99 = trapToDebug ? {{1'd0}, reg_mstatus_spp} : _GEN_80; // @[CSR.scala 671:24]
  assign _GEN_101 = trapToDebug ? reg_mepc : _GEN_83; // @[CSR.scala 671:24]
  assign _GEN_104 = trapToDebug ? reg_mstatus_mpie : _GEN_86; // @[CSR.scala 671:24]
  assign _GEN_105 = trapToDebug ? reg_mstatus_mpp : _GEN_87; // @[CSR.scala 671:24]
  assign _GEN_106 = trapToDebug ? reg_mstatus_mie : _GEN_88; // @[CSR.scala 671:24]
  assign _GEN_108 = exception ? _GEN_90 : reg_dpc; // @[CSR.scala 670:20]
  assign _GEN_112 = exception ? _GEN_94 : reg_sepc; // @[CSR.scala 670:20]
  assign _GEN_116 = exception ? _GEN_98 : reg_mstatus_spie; // @[CSR.scala 670:20]
  assign _GEN_117 = exception ? _GEN_99 : {{1'd0}, reg_mstatus_spp}; // @[CSR.scala 670:20]
  assign _GEN_119 = exception ? _GEN_101 : reg_mepc; // @[CSR.scala 670:20]
  assign _GEN_122 = exception ? _GEN_104 : reg_mstatus_mpie; // @[CSR.scala 670:20]
  assign _GEN_123 = exception ? _GEN_105 : reg_mstatus_mpp; // @[CSR.scala 670:20]
  assign _GEN_124 = exception ? _GEN_106 : reg_mstatus_mie; // @[CSR.scala 670:20]
  assign _GEN_127 = io_rw_addr[10] ? ~_T_650 : ~_T_624; // @[CSR.scala 725:53]
  assign _GEN_132 = ~io_rw_addr[9] | _GEN_116; // @[CSR.scala 719:44]
  assign _GEN_133 = io_rw_addr[9] ? _GEN_117 : 2'h0; // @[CSR.scala 719:44]
  assign _GEN_135 = io_rw_addr[9] ? _GEN_127 : ~_T_857; // @[CSR.scala 719:44]
  assign _GEN_142 = insn_ret ? _GEN_133 : _GEN_117; // @[CSR.scala 718:19]
  assign _T_1942 = _T_980 ? _T_615 : 64'h0; // @[Mux.scala 19:72]
  assign _T_1943 = _T_981 ? _T_620 : 64'h0; // @[Mux.scala 19:72]
  assign _T_1944 = _T_982 ? reg_misa : 64'h0; // @[Mux.scala 19:72]
  assign _T_1945 = _T_983 ? read_mstatus : 64'h0; // @[Mux.scala 19:72]
  assign _T_1946 = _T_984 ? reg_mtvec : 32'h0; // @[Mux.scala 19:72]
  assign _T_1947 = _T_985 ? read_mip : 16'h0; // @[Mux.scala 19:72]
  assign _T_1948 = _T_986 ? reg_mie : 64'h0; // @[Mux.scala 19:72]
  assign _T_1949 = _T_987 ? reg_mscratch : 64'h0; // @[Mux.scala 19:72]
  assign _T_1950 = _T_988 ? _T_629 : 64'h0; // @[Mux.scala 19:72]
  assign _T_1951 = _T_989 ? _T_633 : 64'h0; // @[Mux.scala 19:72]
  assign _T_1952 = _T_990 ? reg_mcause : 64'h0; // @[Mux.scala 19:72]
  assign _T_1953 = _T_991 ? io_hartid : 2'h0; // @[Mux.scala 19:72]
  assign _T_1954 = _T_992 ? _T_646 : 32'h0; // @[Mux.scala 19:72]
  assign _T_1955 = _T_993 ? _T_655 : 64'h0; // @[Mux.scala 19:72]
  assign _T_1956 = _T_994 ? reg_dscratch : 64'h0; // @[Mux.scala 19:72]
  assign _T_1957 = _T_995 ? reg_fflags : 5'h0; // @[Mux.scala 19:72]
  assign _T_1958 = _T_996 ? reg_frm : 3'h0; // @[Mux.scala 19:72]
  assign _T_1959 = _T_997 ? _T_656 : 8'h0; // @[Mux.scala 19:72]
  assign _T_1960 = _T_998 ? _T_303 : 64'h0; // @[Mux.scala 19:72]
  assign _T_1961 = _T_999 ? _T_293 : 64'h0; // @[Mux.scala 19:72]
  assign _T_2049 = _T_1087 ? reg_mcounteren : 32'h0; // @[Mux.scala 19:72]
  assign _T_2050 = _T_1088 ? _T_303 : 64'h0; // @[Mux.scala 19:72]
  assign _T_2051 = _T_1089 ? _T_293 : 64'h0; // @[Mux.scala 19:72]
  assign _T_2052 = _T_1090 ? vpoffset_reg : 27'h0; // @[Mux.scala 19:72]
  assign _T_2053 = _T_1091 ? _T_771 : 32'h0; // @[Mux.scala 19:72]
  assign _T_2054 = _T_1092 ? _T_774 : 32'h0; // @[Mux.scala 19:72]
  assign _T_2055 = _T_1093 ? _T_777 : 32'h0; // @[Mux.scala 19:72]
  assign _T_2056 = _T_1094 ? _T_780 : 32'h0; // @[Mux.scala 19:72]
  assign _T_2057 = _T_1095 ? _T_846[63:0] : 64'h0; // @[Mux.scala 19:72]
  assign _T_2058 = _T_1096 ? _T_782 : 64'h0; // @[Mux.scala 19:72]
  assign _T_2059 = _T_1097 ? _T_781 : 64'h0; // @[Mux.scala 19:72]
  assign _T_2060 = _T_1098 ? reg_sscratch : 64'h0; // @[Mux.scala 19:72]
  assign _T_2061 = _T_1099 ? reg_scause : 64'h0; // @[Mux.scala 19:72]
  assign _T_2062 = _T_1100 ? _T_851 : 64'h0; // @[Mux.scala 19:72]
  assign _T_2063 = _T_1101 ? _T_853 : 64'h0; // @[Mux.scala 19:72]
  assign _T_2064 = _T_1102 ? _T_862 : 64'h0; // @[Mux.scala 19:72]
  assign _T_2065 = _T_1103 ? _T_866 : 64'h0; // @[Mux.scala 19:72]
  assign _T_2066 = _T_1104 ? reg_scounteren : 32'h0; // @[Mux.scala 19:72]
  assign _T_2067 = _T_1105 ? reg_mideleg : 64'h0; // @[Mux.scala 19:72]
  assign _T_2068 = _T_1106 ? reg_medeleg : 64'h0; // @[Mux.scala 19:72]
  assign _T_2069 = _T_1107 ? _T_927 : 64'h0; // @[Mux.scala 19:72]
  assign _T_2071 = _T_1109 ? reg_pmp_0_addr : 30'h0; // @[Mux.scala 19:72]
  assign _T_2072 = _T_1110 ? reg_pmp_1_addr : 30'h0; // @[Mux.scala 19:72]
  assign _T_2073 = _T_1111 ? reg_pmp_2_addr : 30'h0; // @[Mux.scala 19:72]
  assign _T_2074 = _T_1112 ? reg_pmp_3_addr : 30'h0; // @[Mux.scala 19:72]
  assign _T_2075 = _T_1113 ? reg_pmp_4_addr : 30'h0; // @[Mux.scala 19:72]
  assign _T_2076 = _T_1114 ? reg_pmp_5_addr : 30'h0; // @[Mux.scala 19:72]
  assign _T_2077 = _T_1115 ? reg_pmp_6_addr : 30'h0; // @[Mux.scala 19:72]
  assign _T_2078 = _T_1116 ? reg_pmp_7_addr : 30'h0; // @[Mux.scala 19:72]
  assign _T_2088 = _T_1126 ? 64'h1 : 64'h0; // @[Mux.scala 19:72]
  assign _T_2092 = _T_1942 | _T_1943; // @[Mux.scala 19:72]
  assign _T_2093 = _T_2092 | _T_1944; // @[Mux.scala 19:72]
  assign _T_2094 = _T_2093 | _T_1945; // @[Mux.scala 19:72]
  assign _GEN_743 = {{32'd0}, _T_1946}; // @[Mux.scala 19:72]
  assign _T_2095 = _T_2094 | _GEN_743; // @[Mux.scala 19:72]
  assign _GEN_744 = {{48'd0}, _T_1947}; // @[Mux.scala 19:72]
  assign _T_2096 = _T_2095 | _GEN_744; // @[Mux.scala 19:72]
  assign _T_2097 = _T_2096 | _T_1948; // @[Mux.scala 19:72]
  assign _T_2098 = _T_2097 | _T_1949; // @[Mux.scala 19:72]
  assign _T_2099 = _T_2098 | _T_1950; // @[Mux.scala 19:72]
  assign _T_2100 = _T_2099 | _T_1951; // @[Mux.scala 19:72]
  assign _T_2101 = _T_2100 | _T_1952; // @[Mux.scala 19:72]
  assign _GEN_745 = {{62'd0}, _T_1953}; // @[Mux.scala 19:72]
  assign _T_2102 = _T_2101 | _GEN_745; // @[Mux.scala 19:72]
  assign _GEN_746 = {{32'd0}, _T_1954}; // @[Mux.scala 19:72]
  assign _T_2103 = _T_2102 | _GEN_746; // @[Mux.scala 19:72]
  assign _T_2104 = _T_2103 | _T_1955; // @[Mux.scala 19:72]
  assign _T_2105 = _T_2104 | _T_1956; // @[Mux.scala 19:72]
  assign _GEN_747 = {{59'd0}, _T_1957}; // @[Mux.scala 19:72]
  assign _T_2106 = _T_2105 | _GEN_747; // @[Mux.scala 19:72]
  assign _GEN_748 = {{61'd0}, _T_1958}; // @[Mux.scala 19:72]
  assign _T_2107 = _T_2106 | _GEN_748; // @[Mux.scala 19:72]
  assign _GEN_749 = {{56'd0}, _T_1959}; // @[Mux.scala 19:72]
  assign _T_2108 = _T_2107 | _GEN_749; // @[Mux.scala 19:72]
  assign _T_2109 = _T_2108 | _T_1960; // @[Mux.scala 19:72]
  assign _T_2110 = _T_2109 | _T_1961; // @[Mux.scala 19:72]
  assign _GEN_750 = {{32'd0}, _T_2049}; // @[Mux.scala 19:72]
  assign _T_2198 = _T_2110 | _GEN_750; // @[Mux.scala 19:72]
  assign _T_2199 = _T_2198 | _T_2050; // @[Mux.scala 19:72]
  assign _T_2200 = _T_2199 | _T_2051; // @[Mux.scala 19:72]
  assign _GEN_751 = {{37'd0}, _T_2052}; // @[Mux.scala 19:72]
  assign _T_2201 = _T_2200 | _GEN_751; // @[Mux.scala 19:72]
  assign _GEN_752 = {{32'd0}, _T_2053}; // @[Mux.scala 19:72]
  assign _T_2202 = _T_2201 | _GEN_752; // @[Mux.scala 19:72]
  assign _GEN_753 = {{32'd0}, _T_2054}; // @[Mux.scala 19:72]
  assign _T_2203 = _T_2202 | _GEN_753; // @[Mux.scala 19:72]
  assign _GEN_754 = {{32'd0}, _T_2055}; // @[Mux.scala 19:72]
  assign _T_2204 = _T_2203 | _GEN_754; // @[Mux.scala 19:72]
  assign _GEN_755 = {{32'd0}, _T_2056}; // @[Mux.scala 19:72]
  assign _T_2205 = _T_2204 | _GEN_755; // @[Mux.scala 19:72]
  assign _T_2206 = _T_2205 | _T_2057; // @[Mux.scala 19:72]
  assign _T_2207 = _T_2206 | _T_2058; // @[Mux.scala 19:72]
  assign _T_2208 = _T_2207 | _T_2059; // @[Mux.scala 19:72]
  assign _T_2209 = _T_2208 | _T_2060; // @[Mux.scala 19:72]
  assign _T_2210 = _T_2209 | _T_2061; // @[Mux.scala 19:72]
  assign _T_2211 = _T_2210 | _T_2062; // @[Mux.scala 19:72]
  assign _T_2212 = _T_2211 | _T_2063; // @[Mux.scala 19:72]
  assign _T_2213 = _T_2212 | _T_2064; // @[Mux.scala 19:72]
  assign _T_2214 = _T_2213 | _T_2065; // @[Mux.scala 19:72]
  assign _GEN_756 = {{32'd0}, _T_2066}; // @[Mux.scala 19:72]
  assign _T_2215 = _T_2214 | _GEN_756; // @[Mux.scala 19:72]
  assign _T_2216 = _T_2215 | _T_2067; // @[Mux.scala 19:72]
  assign _T_2217 = _T_2216 | _T_2068; // @[Mux.scala 19:72]
  assign _T_2218 = _T_2217 | _T_2069; // @[Mux.scala 19:72]
  assign _GEN_757 = {{34'd0}, _T_2071}; // @[Mux.scala 19:72]
  assign _T_2220 = _T_2218 | _GEN_757; // @[Mux.scala 19:72]
  assign _GEN_758 = {{34'd0}, _T_2072}; // @[Mux.scala 19:72]
  assign _T_2221 = _T_2220 | _GEN_758; // @[Mux.scala 19:72]
  assign _GEN_759 = {{34'd0}, _T_2073}; // @[Mux.scala 19:72]
  assign _T_2222 = _T_2221 | _GEN_759; // @[Mux.scala 19:72]
  assign _GEN_760 = {{34'd0}, _T_2074}; // @[Mux.scala 19:72]
  assign _T_2223 = _T_2222 | _GEN_760; // @[Mux.scala 19:72]
  assign _GEN_761 = {{34'd0}, _T_2075}; // @[Mux.scala 19:72]
  assign _T_2224 = _T_2223 | _GEN_761; // @[Mux.scala 19:72]
  assign _GEN_762 = {{34'd0}, _T_2076}; // @[Mux.scala 19:72]
  assign _T_2225 = _T_2224 | _GEN_762; // @[Mux.scala 19:72]
  assign _GEN_763 = {{34'd0}, _T_2077}; // @[Mux.scala 19:72]
  assign _T_2226 = _T_2225 | _GEN_763; // @[Mux.scala 19:72]
  assign _GEN_764 = {{34'd0}, _T_2078}; // @[Mux.scala 19:72]
  assign _T_2227 = _T_2226 | _GEN_764; // @[Mux.scala 19:72]
  assign _T_2242 = io_rw_cmd == 3'h5; // @[package.scala 14:47]
  assign _T_2243 = io_rw_cmd == 3'h6; // @[package.scala 14:47]
  assign _T_2244 = io_rw_cmd == 3'h7; // @[package.scala 14:47]
  assign _T_3593 = reg_fflags | io_fcsr_flags_bits; // @[CSR.scala 764:30]
  assign _GEN_149 = io_fcsr_flags_valid ? _T_3593 : reg_fflags; // @[CSR.scala 763:30]
  assign _T_3597 = _T_2243 | _T_2244; // @[package.scala 14:62]
  assign csr_wen = _T_3597 | _T_2242; // @[package.scala 14:62]
  assign _GEN_175 = pcode_regs_0_locked ? {{7'd0}, pcode_update_bits_id} : 9'h0; // @[CSR.scala 796:34]
  assign _GEN_176 = pcode_regs_0_locked ? pcode_update_bits_value_base : wdata[31:12]; // @[CSR.scala 796:34]
  assign _GEN_177 = pcode_regs_0_locked ? pcode_update_bits_value_mask : wdata[11:2]; // @[CSR.scala 796:34]
  assign _GEN_178 = pcode_regs_0_locked ? pcode_update_bits_value_valid : wdata[1]; // @[CSR.scala 796:34]
  assign _GEN_179 = pcode_regs_0_locked ? pcode_update_bits_value_locked : wdata[0]; // @[CSR.scala 796:34]
  assign _GEN_184 = _T_1091 & ~pcode_regs_0_locked; // @[CSR.scala 792:40]
  assign _GEN_185 = _T_1091 ? _GEN_175 : {{7'd0}, pcode_update_bits_id}; // @[CSR.scala 792:40]
  assign _GEN_186 = _T_1091 ? _GEN_176 : pcode_update_bits_value_base; // @[CSR.scala 792:40]
  assign _GEN_187 = _T_1091 ? _GEN_177 : pcode_update_bits_value_mask; // @[CSR.scala 792:40]
  assign _GEN_188 = _T_1091 ? _GEN_178 : pcode_update_bits_value_valid; // @[CSR.scala 792:40]
  assign _GEN_189 = _T_1091 ? _GEN_179 : pcode_update_bits_value_locked; // @[CSR.scala 792:40]
  assign _GEN_214 = ~pcode_regs_1_locked | _GEN_184; // @[CSR.scala 796:34]
  assign _GEN_215 = pcode_regs_1_locked ? _GEN_185 : 9'h1; // @[CSR.scala 796:34]
  assign _GEN_224 = _T_1092 ? _GEN_214 : _GEN_184; // @[CSR.scala 792:40]
  assign _GEN_225 = _T_1092 ? _GEN_215 : _GEN_185; // @[CSR.scala 792:40]
  assign _GEN_254 = ~pcode_regs_2_locked | _GEN_224; // @[CSR.scala 796:34]
  assign _GEN_255 = pcode_regs_2_locked ? _GEN_225 : 9'h2; // @[CSR.scala 796:34]
  assign _GEN_264 = _T_1093 ? _GEN_254 : _GEN_224; // @[CSR.scala 792:40]
  assign _GEN_265 = _T_1093 ? _GEN_255 : _GEN_225; // @[CSR.scala 792:40]
  assign _GEN_294 = ~pcode_regs_3_locked | _GEN_264; // @[CSR.scala 796:34]
  assign _GEN_295 = pcode_regs_3_locked ? _GEN_265 : 9'h3; // @[CSR.scala 796:34]
  assign _GEN_304 = _T_1094 ? _GEN_294 : _GEN_264; // @[CSR.scala 792:40]
  assign _GEN_305 = _T_1094 ? _GEN_295 : _GEN_265; // @[CSR.scala 792:40]
  assign _T_3676 = {{37'd0}, wdata};
  assign _T_3706 = _T_3676[12:11] == 2'h2; // @[CSR.scala 1035:27]
  assign _T_3708 = _T_3676[14:13] != 2'h0; // @[CSR.scala 1055:73]
  assign _GEN_320 = _T_983 ? {{1'd0}, _T_3676[8]} : _GEN_142; // @[CSR.scala 814:39]
  assign _T_3716 = ~io_pc[1] | wdata[2]; // @[CSR.scala 841:43]
  assign _T_3719 = {~wdata[5], 3'h0}; // @[CSR.scala 843:38]
  assign _GEN_765 = {{60'd0}, _T_3719}; // @[CSR.scala 843:32]
  assign _T_3720 = ~wdata | _GEN_765; // @[CSR.scala 843:32]
  assign _T_3722 = ~_T_3720 & 64'h102d; // @[CSR.scala 843:55]
  assign _T_3724 = reg_misa & 64'hffffffffffffefd2; // @[CSR.scala 843:73]
  assign _T_3725 = _T_3722 | _T_3724; // @[CSR.scala 843:62]
  assign _T_3740 = {4'h0,2'h0,reg_mip_seip,1'h0,2'h0,reg_mip_stip,1'h0,2'h0,reg_mip_ssip,1'h0}; // @[CSR.scala 851:59]
  assign _T_3742 = io_rw_cmd[1] ? _T_3740 : 16'h0; // @[CSR.scala 1031:9]
  assign _GEN_766 = {{48'd0}, _T_3742}; // @[CSR.scala 1031:34]
  assign _T_3743 = _GEN_766 | io_rw_wdata; // @[CSR.scala 1031:34]
  assign _T_3749 = _T_3743 & ~_T_1135; // @[CSR.scala 1031:43]
  assign _T_3777 = wdata & 64'haaa; // @[CSR.scala 858:59]
  assign _T_3779 = ~wdata | 64'h1; // @[CSR.scala 1052:31]
  assign _GEN_333 = _T_988 ? ~_T_3779 : {{24'd0}, _GEN_119}; // @[CSR.scala 859:40]
  assign _T_3782 = ~wdata | 64'h2; // @[CSR.scala 862:64]
  assign _T_3784 = wdata[0] ? 8'hfc : 8'h0; // @[CSR.scala 862:75]
  assign _GEN_767 = {{56'd0}, _T_3784}; // @[CSR.scala 862:70]
  assign _T_3785 = _T_3782 | _GEN_767; // @[CSR.scala 862:70]
  assign _GEN_335 = _T_984 ? ~_T_3785 : {{32'd0}, reg_mtvec}; // @[CSR.scala 862:40]
  assign _T_3787 = wdata & 64'h800000000000000f; // @[CSR.scala 863:62]
  assign _GEN_338 = _T_998 ? wdata : {{57'd0}, _T_297}; // @[CSR.scala 1049:31]
  assign _GEN_340 = _T_999 ? wdata : {{57'd0}, _T_287}; // @[CSR.scala 1049:31]
  assign _GEN_343 = _T_995 ? wdata : {{59'd0}, _GEN_149}; // @[CSR.scala 876:40]
  assign _GEN_345 = _T_996 ? wdata : {{61'd0}, reg_frm}; // @[CSR.scala 877:40]
  assign _GEN_347 = _T_997 ? wdata : _GEN_343; // @[CSR.scala 878:40]
  assign _GEN_348 = _T_997 ? {{5'd0}, wdata[63:5]} : _GEN_345; // @[CSR.scala 878:40]
  assign _T_3813 = wdata[1:0] == 2'h2; // @[CSR.scala 1035:27]
  assign _GEN_354 = _T_993 ? ~_T_3779 : {{24'd0}, _GEN_108}; // @[CSR.scala 889:42]
  assign _GEN_358 = _T_1095 ? {{1'd0}, _T_3676[8]} : _GEN_320; // @[CSR.scala 893:41]
  assign _T_3859 = _GEN_730 & ~reg_mideleg; // @[CSR.scala 904:52]
  assign _T_3860 = wdata & reg_mideleg; // @[CSR.scala 904:77]
  assign _T_3861 = _T_3859 | _T_3860; // @[CSR.scala 904:68]
  assign _T_3894 = wdata[63:60] == 4'h0; // @[CSR.scala 910:30]
  assign _T_3895 = wdata[63:60] == 4'h8; // @[CSR.scala 911:30]
  assign _T_3898 = _T_3894 | _T_3895; // @[CSR.scala 912:36]
  assign _T_3901 = reg_mie & ~reg_mideleg; // @[CSR.scala 917:64]
  assign _T_3903 = _T_3901 | _T_3860; // @[CSR.scala 917:80]
  assign _GEN_370 = _T_1102 ? ~_T_3779 : {{24'd0}, _GEN_112}; // @[CSR.scala 919:42]
  assign _GEN_371 = _T_1103 ? ~_T_3785 : {{25'd0}, reg_stvec}; // @[CSR.scala 920:42]
  assign _T_3913 = wdata & 64'h800000000000001f; // @[CSR.scala 921:64]
  assign _T_3915 = wdata & 64'h222; // @[CSR.scala 923:65]
  assign _T_3916 = wdata & 64'hb109; // @[CSR.scala 924:65]
  assign _T_3917 = wdata & 64'h7; // @[CSR.scala 925:70]
  assign _GEN_376 = _T_1104 ? _T_3917 : {{32'd0}, reg_scounteren}; // @[CSR.scala 925:44]
  assign _GEN_377 = _T_1087 ? _T_3917 : {{32'd0}, reg_mcounteren}; // @[CSR.scala 928:44]
  assign _T_3921 = ~reg_bp_0_control_dmode | reg_debug; // @[CSR.scala 934:31]
  assign _T_3942 = wdata[59] & reg_debug; // @[CSR.scala 937:36]
  assign _T_3943 = _T_3942 & wdata[12]; // @[CSR.scala 940:38]
  assign _T_3945 = _T_1107 & ~reg_pmp_0_cfg_l; // @[CSR.scala 947:57]
  assign _T_3961 = ~reg_pmp_1_cfg_a[1] & reg_pmp_1_cfg_a[0]; // @[PMP.scala 41:20]
  assign _T_3962 = reg_pmp_1_cfg_l & _T_3961; // @[PMP.scala 43:62]
  assign _T_3963 = reg_pmp_0_cfg_l | _T_3962; // @[PMP.scala 43:44]
  assign _T_3965 = _T_1109 & ~_T_3963; // @[CSR.scala 954:45]
  assign _GEN_485 = _T_3965 ? wdata : {{34'd0}, reg_pmp_0_addr}; // @[CSR.scala 954:71]
  assign _T_3967 = _T_1107 & ~reg_pmp_1_cfg_l; // @[CSR.scala 947:57]
  assign _T_3983 = ~reg_pmp_2_cfg_a[1] & reg_pmp_2_cfg_a[0]; // @[PMP.scala 41:20]
  assign _T_3984 = reg_pmp_2_cfg_l & _T_3983; // @[PMP.scala 43:62]
  assign _T_3985 = reg_pmp_1_cfg_l | _T_3984; // @[PMP.scala 43:44]
  assign _T_3987 = _T_1110 & ~_T_3985; // @[CSR.scala 954:45]
  assign _GEN_492 = _T_3987 ? wdata : {{34'd0}, reg_pmp_1_addr}; // @[CSR.scala 954:71]
  assign _T_3989 = _T_1107 & ~reg_pmp_2_cfg_l; // @[CSR.scala 947:57]
  assign _T_4005 = ~reg_pmp_3_cfg_a[1] & reg_pmp_3_cfg_a[0]; // @[PMP.scala 41:20]
  assign _T_4006 = reg_pmp_3_cfg_l & _T_4005; // @[PMP.scala 43:62]
  assign _T_4007 = reg_pmp_2_cfg_l | _T_4006; // @[PMP.scala 43:44]
  assign _T_4009 = _T_1111 & ~_T_4007; // @[CSR.scala 954:45]
  assign _GEN_499 = _T_4009 ? wdata : {{34'd0}, reg_pmp_2_addr}; // @[CSR.scala 954:71]
  assign _T_4011 = _T_1107 & ~reg_pmp_3_cfg_l; // @[CSR.scala 947:57]
  assign _T_4027 = ~reg_pmp_4_cfg_a[1] & reg_pmp_4_cfg_a[0]; // @[PMP.scala 41:20]
  assign _T_4028 = reg_pmp_4_cfg_l & _T_4027; // @[PMP.scala 43:62]
  assign _T_4029 = reg_pmp_3_cfg_l | _T_4028; // @[PMP.scala 43:44]
  assign _T_4031 = _T_1112 & ~_T_4029; // @[CSR.scala 954:45]
  assign _GEN_506 = _T_4031 ? wdata : {{34'd0}, reg_pmp_3_addr}; // @[CSR.scala 954:71]
  assign _T_4033 = _T_1107 & ~reg_pmp_4_cfg_l; // @[CSR.scala 947:57]
  assign _T_4049 = ~reg_pmp_5_cfg_a[1] & reg_pmp_5_cfg_a[0]; // @[PMP.scala 41:20]
  assign _T_4050 = reg_pmp_5_cfg_l & _T_4049; // @[PMP.scala 43:62]
  assign _T_4051 = reg_pmp_4_cfg_l | _T_4050; // @[PMP.scala 43:44]
  assign _T_4053 = _T_1113 & ~_T_4051; // @[CSR.scala 954:45]
  assign _GEN_513 = _T_4053 ? wdata : {{34'd0}, reg_pmp_4_addr}; // @[CSR.scala 954:71]
  assign _T_4055 = _T_1107 & ~reg_pmp_5_cfg_l; // @[CSR.scala 947:57]
  assign _T_4071 = ~reg_pmp_6_cfg_a[1] & reg_pmp_6_cfg_a[0]; // @[PMP.scala 41:20]
  assign _T_4072 = reg_pmp_6_cfg_l & _T_4071; // @[PMP.scala 43:62]
  assign _T_4073 = reg_pmp_5_cfg_l | _T_4072; // @[PMP.scala 43:44]
  assign _T_4075 = _T_1114 & ~_T_4073; // @[CSR.scala 954:45]
  assign _GEN_520 = _T_4075 ? wdata : {{34'd0}, reg_pmp_5_addr}; // @[CSR.scala 954:71]
  assign _T_4077 = _T_1107 & ~reg_pmp_6_cfg_l; // @[CSR.scala 947:57]
  assign _T_4093 = ~reg_pmp_7_cfg_a[1] & reg_pmp_7_cfg_a[0]; // @[PMP.scala 41:20]
  assign _T_4094 = reg_pmp_7_cfg_l & _T_4093; // @[PMP.scala 43:62]
  assign _T_4095 = reg_pmp_6_cfg_l | _T_4094; // @[PMP.scala 43:44]
  assign _T_4097 = _T_1115 & ~_T_4095; // @[CSR.scala 954:45]
  assign _GEN_527 = _T_4097 ? wdata : {{34'd0}, reg_pmp_6_addr}; // @[CSR.scala 954:71]
  assign _T_4099 = _T_1107 & ~reg_pmp_7_cfg_l; // @[CSR.scala 947:57]
  assign _T_4117 = reg_pmp_7_cfg_l | _T_4094; // @[PMP.scala 43:44]
  assign _T_4119 = _T_1116 & ~_T_4117; // @[CSR.scala 954:45]
  assign _GEN_534 = _T_4119 ? wdata : {{34'd0}, reg_pmp_7_addr}; // @[CSR.scala 954:71]
  assign _GEN_547 = csr_wen ? _GEN_305 : {{7'd0}, pcode_update_bits_id}; // @[CSR.scala 782:18]
  assign _GEN_562 = csr_wen ? _GEN_358 : _GEN_142; // @[CSR.scala 782:18]
  assign _GEN_574 = csr_wen ? _GEN_333 : {{24'd0}, _GEN_119}; // @[CSR.scala 782:18]
  assign _GEN_576 = csr_wen ? _GEN_335 : {{32'd0}, reg_mtvec}; // @[CSR.scala 782:18]
  assign _GEN_579 = csr_wen ? _GEN_338 : {{57'd0}, _T_297}; // @[CSR.scala 782:18]
  assign _GEN_581 = csr_wen ? _GEN_340 : {{57'd0}, _T_287}; // @[CSR.scala 782:18]
  assign _GEN_584 = csr_wen ? _GEN_347 : {{59'd0}, _GEN_149}; // @[CSR.scala 782:18]
  assign _GEN_585 = csr_wen ? _GEN_348 : {{61'd0}, reg_frm}; // @[CSR.scala 782:18]
  assign _GEN_591 = csr_wen ? _GEN_354 : {{24'd0}, _GEN_108}; // @[CSR.scala 782:18]
  assign _GEN_596 = csr_wen ? _GEN_370 : {{24'd0}, _GEN_112}; // @[CSR.scala 782:18]
  assign _GEN_597 = csr_wen ? _GEN_371 : {{25'd0}, reg_stvec}; // @[CSR.scala 782:18]
  assign _GEN_602 = csr_wen ? _GEN_376 : {{32'd0}, reg_scounteren}; // @[CSR.scala 782:18]
  assign _GEN_603 = csr_wen ? _GEN_377 : {{32'd0}, reg_mcounteren}; // @[CSR.scala 782:18]
  assign _GEN_643 = csr_wen ? _GEN_485 : {{34'd0}, reg_pmp_0_addr}; // @[CSR.scala 782:18]
  assign _GEN_650 = csr_wen ? _GEN_492 : {{34'd0}, reg_pmp_1_addr}; // @[CSR.scala 782:18]
  assign _GEN_657 = csr_wen ? _GEN_499 : {{34'd0}, reg_pmp_2_addr}; // @[CSR.scala 782:18]
  assign _GEN_664 = csr_wen ? _GEN_506 : {{34'd0}, reg_pmp_3_addr}; // @[CSR.scala 782:18]
  assign _GEN_671 = csr_wen ? _GEN_513 : {{34'd0}, reg_pmp_4_addr}; // @[CSR.scala 782:18]
  assign _GEN_678 = csr_wen ? _GEN_520 : {{34'd0}, reg_pmp_5_addr}; // @[CSR.scala 782:18]
  assign _GEN_685 = csr_wen ? _GEN_527 : {{34'd0}, reg_pmp_6_addr}; // @[CSR.scala 782:18]
  assign _GEN_692 = csr_wen ? _GEN_534 : {{34'd0}, reg_pmp_7_addr}; // @[CSR.scala 782:18]
  assign io_rw_rdata = _T_2227 | _T_2088; // @[CSR.scala 747:15]
  assign io_pcode_req_valid = pcode_update_valid; // @[CSR.scala 502:18]
  assign io_pcode_req_bits_id = pcode_update_bits_id; // @[CSR.scala 502:18]
  assign io_pcode_req_bits_value_base = pcode_update_bits_value_base; // @[CSR.scala 502:18]
  assign io_pcode_req_bits_value_mask = pcode_update_bits_value_mask; // @[CSR.scala 502:18]
  assign io_pcode_req_bits_value_valid = pcode_update_bits_value_valid; // @[CSR.scala 502:18]
  assign io_pcode_req_bits_value_locked = pcode_update_bits_value_locked; // @[CSR.scala 502:18]
  assign io_vpoffset_req_bits_value = vpoffset_update_bits_value; // @[CSR.scala 498:21]
  assign io_decode_0_fp_illegal = _T_1208 | ~reg_misa[5]; // @[CSR.scala 601:23]
  assign io_decode_0_fp_csr = _T_1212 == 12'h0; // @[CSR.scala 602:19]
  assign io_decode_0_read_illegal = _T_1546 | _T_1547; // @[CSR.scala 604:25]
  assign io_decode_0_write_illegal = ~io_decode_0_csr[11:10] == 2'h0; // @[CSR.scala 610:26]
  assign io_decode_0_write_flush = ~_T_1558; // @[CSR.scala 611:24]
  assign io_decode_0_system_illegal = _T_1567 | _T_1569; // @[CSR.scala 612:27]
  assign io_csr_stall = reg_wfi; // @[CSR.scala 739:16]
  assign io_eret = _T_1627 | insn_ret; // @[CSR.scala 643:11]
  assign io_singleStep = reg_dcsr_step & ~reg_debug; // @[CSR.scala 644:17]
  assign io_status_debug = reg_debug; // @[CSR.scala 645:13 CSR.scala 647:19]
  assign io_status_isa = reg_misa[31:0]; // @[CSR.scala 645:13 CSR.scala 648:17]
  assign io_status_dprv = _T_1626; // @[CSR.scala 645:13 CSR.scala 651:18]
  assign io_status_prv = reg_mstatus_prv; // @[CSR.scala 645:13]
  assign io_status_sd = _T_1618 | _T_1620; // @[CSR.scala 645:13 CSR.scala 646:16]
  assign io_status_zero2 = 27'h0; // @[CSR.scala 645:13]
  assign io_status_sxl = 2'h2; // @[CSR.scala 645:13 CSR.scala 650:17]
  assign io_status_uxl = 2'h2; // @[CSR.scala 645:13 CSR.scala 649:17]
  assign io_status_sd_rv32 = 1'h0; // @[CSR.scala 645:13]
  assign io_status_zero1 = 8'h0; // @[CSR.scala 645:13]
  assign io_status_tsr = reg_mstatus_tsr; // @[CSR.scala 645:13]
  assign io_status_tw = reg_mstatus_tw; // @[CSR.scala 645:13]
  assign io_status_tvm = reg_mstatus_tvm; // @[CSR.scala 645:13]
  assign io_status_mxr = reg_mstatus_mxr; // @[CSR.scala 645:13]
  assign io_status_sum = reg_mstatus_sum; // @[CSR.scala 645:13]
  assign io_status_mprv = reg_mstatus_mprv; // @[CSR.scala 645:13]
  assign io_status_xs = 2'h0; // @[CSR.scala 645:13]
  assign io_status_fs = reg_mstatus_fs; // @[CSR.scala 645:13]
  assign io_status_mpp = reg_mstatus_mpp; // @[CSR.scala 645:13]
  assign io_status_hpp = 2'h0; // @[CSR.scala 645:13]
  assign io_status_spp = reg_mstatus_spp; // @[CSR.scala 645:13]
  assign io_status_mpie = reg_mstatus_mpie; // @[CSR.scala 645:13]
  assign io_status_hpie = 1'h0; // @[CSR.scala 645:13]
  assign io_status_spie = reg_mstatus_spie; // @[CSR.scala 645:13]
  assign io_status_upie = 1'h0; // @[CSR.scala 645:13]
  assign io_status_mie = reg_mstatus_mie; // @[CSR.scala 645:13]
  assign io_status_hie = 1'h0; // @[CSR.scala 645:13]
  assign io_status_sie = reg_mstatus_sie; // @[CSR.scala 645:13]
  assign io_status_uie = 1'h0; // @[CSR.scala 645:13]
  assign io_ptbr_mode = reg_sptbr_mode; // @[CSR.scala 642:11]
  assign io_ptbr_ppn = reg_sptbr_ppn; // @[CSR.scala 642:11]
  assign io_evec = insn_ret ? _GEN_135 : tvec; // @[CSR.scala 641:11 CSR.scala 724:15 CSR.scala 728:15 CSR.scala 734:15]
  assign io_fcsr_rm = reg_frm; // @[CSR.scala 762:14]
  assign io_interrupt = _T_489 & ~reg_debug; // @[CSR.scala 382:16]
  assign io_interrupt_cause = 64'h8000000000000000 + _GEN_731; // @[CSR.scala 383:22]
  assign io_bp_0_control_action = reg_bp_0_control_action; // @[CSR.scala 384:9]
  assign io_bp_0_control_tmatch = reg_bp_0_control_tmatch; // @[CSR.scala 384:9]
  assign io_bp_0_control_m = reg_bp_0_control_m; // @[CSR.scala 384:9]
  assign io_bp_0_control_s = reg_bp_0_control_s; // @[CSR.scala 384:9]
  assign io_bp_0_control_u = reg_bp_0_control_u; // @[CSR.scala 384:9]
  assign io_bp_0_control_x = reg_bp_0_control_x; // @[CSR.scala 384:9]
  assign io_bp_0_control_w = reg_bp_0_control_w; // @[CSR.scala 384:9]
  assign io_bp_0_control_r = reg_bp_0_control_r; // @[CSR.scala 384:9]
  assign io_bp_0_address = reg_bp_0_address; // @[CSR.scala 384:9]
  assign io_pmp_0_cfg_l = reg_pmp_0_cfg_l; // @[CSR.scala 385:10]
  assign io_pmp_0_cfg_a = reg_pmp_0_cfg_a; // @[CSR.scala 385:10]
  assign io_pmp_0_cfg_x = reg_pmp_0_cfg_x; // @[CSR.scala 385:10]
  assign io_pmp_0_cfg_w = reg_pmp_0_cfg_w; // @[CSR.scala 385:10]
  assign io_pmp_0_cfg_r = reg_pmp_0_cfg_r; // @[CSR.scala 385:10]
  assign io_pmp_0_addr = reg_pmp_0_addr; // @[CSR.scala 385:10]
  assign io_pmp_0_mask = _T_501[31:0]; // @[CSR.scala 385:10]
  assign io_pmp_1_cfg_l = reg_pmp_1_cfg_l; // @[CSR.scala 385:10]
  assign io_pmp_1_cfg_a = reg_pmp_1_cfg_a; // @[CSR.scala 385:10]
  assign io_pmp_1_cfg_x = reg_pmp_1_cfg_x; // @[CSR.scala 385:10]
  assign io_pmp_1_cfg_w = reg_pmp_1_cfg_w; // @[CSR.scala 385:10]
  assign io_pmp_1_cfg_r = reg_pmp_1_cfg_r; // @[CSR.scala 385:10]
  assign io_pmp_1_addr = reg_pmp_1_addr; // @[CSR.scala 385:10]
  assign io_pmp_1_mask = _T_511[31:0]; // @[CSR.scala 385:10]
  assign io_pmp_2_cfg_l = reg_pmp_2_cfg_l; // @[CSR.scala 385:10]
  assign io_pmp_2_cfg_a = reg_pmp_2_cfg_a; // @[CSR.scala 385:10]
  assign io_pmp_2_cfg_x = reg_pmp_2_cfg_x; // @[CSR.scala 385:10]
  assign io_pmp_2_cfg_w = reg_pmp_2_cfg_w; // @[CSR.scala 385:10]
  assign io_pmp_2_cfg_r = reg_pmp_2_cfg_r; // @[CSR.scala 385:10]
  assign io_pmp_2_addr = reg_pmp_2_addr; // @[CSR.scala 385:10]
  assign io_pmp_2_mask = _T_521[31:0]; // @[CSR.scala 385:10]
  assign io_pmp_3_cfg_l = reg_pmp_3_cfg_l; // @[CSR.scala 385:10]
  assign io_pmp_3_cfg_a = reg_pmp_3_cfg_a; // @[CSR.scala 385:10]
  assign io_pmp_3_cfg_x = reg_pmp_3_cfg_x; // @[CSR.scala 385:10]
  assign io_pmp_3_cfg_w = reg_pmp_3_cfg_w; // @[CSR.scala 385:10]
  assign io_pmp_3_cfg_r = reg_pmp_3_cfg_r; // @[CSR.scala 385:10]
  assign io_pmp_3_addr = reg_pmp_3_addr; // @[CSR.scala 385:10]
  assign io_pmp_3_mask = _T_531[31:0]; // @[CSR.scala 385:10]
  assign io_pmp_4_cfg_l = reg_pmp_4_cfg_l; // @[CSR.scala 385:10]
  assign io_pmp_4_cfg_a = reg_pmp_4_cfg_a; // @[CSR.scala 385:10]
  assign io_pmp_4_cfg_x = reg_pmp_4_cfg_x; // @[CSR.scala 385:10]
  assign io_pmp_4_cfg_w = reg_pmp_4_cfg_w; // @[CSR.scala 385:10]
  assign io_pmp_4_cfg_r = reg_pmp_4_cfg_r; // @[CSR.scala 385:10]
  assign io_pmp_4_addr = reg_pmp_4_addr; // @[CSR.scala 385:10]
  assign io_pmp_4_mask = _T_541[31:0]; // @[CSR.scala 385:10]
  assign io_pmp_5_cfg_l = reg_pmp_5_cfg_l; // @[CSR.scala 385:10]
  assign io_pmp_5_cfg_a = reg_pmp_5_cfg_a; // @[CSR.scala 385:10]
  assign io_pmp_5_cfg_x = reg_pmp_5_cfg_x; // @[CSR.scala 385:10]
  assign io_pmp_5_cfg_w = reg_pmp_5_cfg_w; // @[CSR.scala 385:10]
  assign io_pmp_5_cfg_r = reg_pmp_5_cfg_r; // @[CSR.scala 385:10]
  assign io_pmp_5_addr = reg_pmp_5_addr; // @[CSR.scala 385:10]
  assign io_pmp_5_mask = _T_551[31:0]; // @[CSR.scala 385:10]
  assign io_pmp_6_cfg_l = reg_pmp_6_cfg_l; // @[CSR.scala 385:10]
  assign io_pmp_6_cfg_a = reg_pmp_6_cfg_a; // @[CSR.scala 385:10]
  assign io_pmp_6_cfg_x = reg_pmp_6_cfg_x; // @[CSR.scala 385:10]
  assign io_pmp_6_cfg_w = reg_pmp_6_cfg_w; // @[CSR.scala 385:10]
  assign io_pmp_6_cfg_r = reg_pmp_6_cfg_r; // @[CSR.scala 385:10]
  assign io_pmp_6_addr = reg_pmp_6_addr; // @[CSR.scala 385:10]
  assign io_pmp_6_mask = _T_561[31:0]; // @[CSR.scala 385:10]
  assign io_pmp_7_cfg_l = reg_pmp_7_cfg_l; // @[CSR.scala 385:10]
  assign io_pmp_7_cfg_a = reg_pmp_7_cfg_a; // @[CSR.scala 385:10]
  assign io_pmp_7_cfg_x = reg_pmp_7_cfg_x; // @[CSR.scala 385:10]
  assign io_pmp_7_cfg_w = reg_pmp_7_cfg_w; // @[CSR.scala 385:10]
  assign io_pmp_7_cfg_r = reg_pmp_7_cfg_r; // @[CSR.scala 385:10]
  assign io_pmp_7_addr = reg_pmp_7_addr; // @[CSR.scala 385:10]
  assign io_pmp_7_mask = _T_571[31:0]; // @[CSR.scala 385:10]
  assign CSRFile_cov_read_addr = CSRFile_state;
  assign CSRFile_cov_read_data = CSRFile_cov[CSRFile_cov_read_addr]; // @[Coverage map for CSRFile]
  assign CSRFile_cov_write_data = 1'h1;
  assign CSRFile_cov_write_addr = CSRFile_state;
  assign CSRFile_cov_write_mask = 1'h1;
  assign CSRFile_cov_write_en = 1'h1;
  assign reg_singleStepped_shl = {reg_singleStepped, 15'h0};
  assign reg_singleStepped_pad = {4'h0,reg_singleStepped_shl};
  assign reg_debug_shl = reg_debug;
  assign reg_debug_pad = {19'h0,reg_debug_shl};
  assign reg_pmp_7_cfg_a_shl = {reg_pmp_7_cfg_a, 8'h0};
  assign reg_pmp_7_cfg_a_pad = {10'h0,reg_pmp_7_cfg_a_shl};
  assign reg_dcsr_ebreaku_shl = {reg_dcsr_ebreaku, 17'h0};
  assign reg_dcsr_ebreaku_pad = {2'h0,reg_dcsr_ebreaku_shl};
  assign reg_dcsr_ebreaks_shl = {reg_dcsr_ebreaks, 13'h0};
  assign reg_dcsr_ebreaks_pad = {6'h0,reg_dcsr_ebreaks_shl};
  assign reg_pmp_6_cfg_l_shl = {reg_pmp_6_cfg_l, 7'h0};
  assign reg_pmp_6_cfg_l_pad = {12'h0,reg_pmp_6_cfg_l_shl};
  assign reg_mstatus_mie_shl = {reg_mstatus_mie, 14'h0};
  assign reg_mstatus_mie_pad = {5'h0,reg_mstatus_mie_shl};
  assign reg_pmp_2_cfg_l_shl = {reg_pmp_2_cfg_l, 7'h0};
  assign reg_pmp_2_cfg_l_pad = {12'h0,reg_pmp_2_cfg_l_shl};
  assign reg_mstatus_mprv_shl = reg_mstatus_mprv;
  assign reg_mstatus_mprv_pad = {19'h0,reg_mstatus_mprv_shl};
  assign reg_pmp_0_cfg_l_shl = {reg_pmp_0_cfg_l, 14'h0};
  assign reg_pmp_0_cfg_l_pad = {5'h0,reg_pmp_0_cfg_l_shl};
  assign _T_310_shl = {_T_310, 7'h0};
  assign _T_310_pad = {12'h0,_T_310_shl};
  assign reg_pmp_3_cfg_l_shl = {reg_pmp_3_cfg_l, 11'h0};
  assign reg_pmp_3_cfg_l_pad = {8'h0,reg_pmp_3_cfg_l_shl};
  assign reg_mip_stip_shl = {reg_mip_stip, 14'h0};
  assign reg_mip_stip_pad = {5'h0,reg_mip_stip_shl};
  assign reg_mip_ssip_shl = reg_mip_ssip;
  assign reg_mip_ssip_pad = {19'h0,reg_mip_ssip_shl};
  assign reg_pmp_5_cfg_l_shl = {reg_pmp_5_cfg_l, 19'h0};
  assign reg_pmp_5_cfg_l_pad = reg_pmp_5_cfg_l_shl;
  assign reg_mstatus_spp_shl = {reg_mstatus_spp, 6'h0};
  assign reg_mstatus_spp_pad = {13'h0,reg_mstatus_spp_shl};
  assign reg_pmp_4_cfg_l_shl = {reg_pmp_4_cfg_l, 3'h0};
  assign reg_pmp_4_cfg_l_pad = {16'h0,reg_pmp_4_cfg_l_shl};
  assign reg_dcsr_ebreakm_shl = {reg_dcsr_ebreakm, 5'h0};
  assign reg_dcsr_ebreakm_pad = {14'h0,reg_dcsr_ebreakm_shl};
  assign reg_mip_seip_shl = {reg_mip_seip, 13'h0};
  assign reg_mip_seip_pad = {6'h0,reg_mip_seip_shl};
  assign reg_pmp_1_cfg_l_shl = {reg_pmp_1_cfg_l, 16'h0};
  assign reg_pmp_1_cfg_l_pad = {3'h0,reg_pmp_1_cfg_l_shl};
  assign reg_bp_0_control_dmode_shl = {reg_bp_0_control_dmode, 11'h0};
  assign reg_bp_0_control_dmode_pad = {8'h0,reg_bp_0_control_dmode_shl};
  assign reg_pmp_7_cfg_l_shl = {reg_pmp_7_cfg_l, 7'h0};
  assign reg_pmp_7_cfg_l_pad = {12'h0,reg_pmp_7_cfg_l_shl};
  assign reg_mstatus_prv_shl = {reg_mstatus_prv, 2'h0};
  assign reg_mstatus_prv_pad = {16'h0,reg_mstatus_prv_shl};
  assign reg_wfi_shl = {reg_wfi, 19'h0};
  assign reg_wfi_pad = reg_wfi_shl;
  assign reg_mstatus_sie_shl = {reg_mstatus_sie, 3'h0};
  assign reg_mstatus_sie_pad = {16'h0,reg_mstatus_sie_shl};
  assign pcode_regs_0_locked_shl = {pcode_regs_0_locked, 15'h0};
  assign pcode_regs_0_locked_pad = {4'h0,pcode_regs_0_locked_shl};
  assign pcode_regs_1_locked_shl = {pcode_regs_1_locked, 15'h0};
  assign pcode_regs_1_locked_pad = {4'h0,pcode_regs_1_locked_shl};
  assign pcode_regs_2_locked_shl = {pcode_regs_2_locked, 15'h0};
  assign pcode_regs_2_locked_pad = {4'h0,pcode_regs_2_locked_shl};
  assign pcode_regs_3_locked_shl = {pcode_regs_3_locked, 15'h0};
  assign pcode_regs_3_locked_pad = {4'h0,pcode_regs_3_locked_shl};
  assign CSRFile_xor16 = reg_debug_pad ^ reg_pmp_7_cfg_a_pad;
  assign CSRFile_xor7 = reg_singleStepped_pad ^ CSRFile_xor16;
  assign CSRFile_xor17 = reg_dcsr_ebreaku_pad ^ reg_dcsr_ebreaks_pad;
  assign CSRFile_xor18 = reg_pmp_6_cfg_l_pad ^ reg_mstatus_mie_pad;
  assign CSRFile_xor8 = CSRFile_xor17 ^ CSRFile_xor18;
  assign CSRFile_xor3 = CSRFile_xor7 ^ CSRFile_xor8;
  assign CSRFile_xor20 = reg_mstatus_mprv_pad ^ reg_pmp_0_cfg_l_pad;
  assign CSRFile_xor9 = reg_pmp_2_cfg_l_pad ^ CSRFile_xor20;
  assign CSRFile_xor21 = _T_310_pad ^ reg_pmp_3_cfg_l_pad;
  assign CSRFile_xor22 = reg_mip_stip_pad ^ reg_mip_ssip_pad;
  assign CSRFile_xor10 = CSRFile_xor21 ^ CSRFile_xor22;
  assign CSRFile_xor4 = CSRFile_xor9 ^ CSRFile_xor10;
  assign CSRFile_xor1 = CSRFile_xor3 ^ CSRFile_xor4;
  assign CSRFile_xor24 = reg_mstatus_spp_pad ^ reg_pmp_4_cfg_l_pad;
  assign CSRFile_xor11 = reg_pmp_5_cfg_l_pad ^ CSRFile_xor24;
  assign CSRFile_xor25 = reg_dcsr_ebreakm_pad ^ reg_mip_seip_pad;
  assign CSRFile_xor26 = reg_pmp_1_cfg_l_pad ^ reg_bp_0_control_dmode_pad;
  assign CSRFile_xor12 = CSRFile_xor25 ^ CSRFile_xor26;
  assign CSRFile_xor5 = CSRFile_xor11 ^ CSRFile_xor12;
  assign CSRFile_xor27 = reg_pmp_7_cfg_l_pad ^ reg_mstatus_prv_pad;
  assign CSRFile_xor28 = reg_wfi_pad ^ reg_mstatus_sie_pad;
  assign CSRFile_xor13 = CSRFile_xor27 ^ CSRFile_xor28;
  assign CSRFile_xor29 = pcode_regs_0_locked_pad ^ pcode_regs_1_locked_pad;
  assign CSRFile_xor30 = pcode_regs_2_locked_pad ^ pcode_regs_3_locked_pad;
  assign CSRFile_xor14 = CSRFile_xor29 ^ CSRFile_xor30;
  assign CSRFile_xor6 = CSRFile_xor13 ^ CSRFile_xor14;
  assign CSRFile_xor2 = CSRFile_xor5 ^ CSRFile_xor6;
  assign CSRFile_xor0 = CSRFile_xor1 ^ CSRFile_xor2;
  assign io_covSum = CSRFile_covSum;
  assign stopEn0 = ~_T_1633;
  assign stopEn1 = ~_T_1655;
  assign CSRFile_or0 = stopEn0 | stopEn1;
  assign metaAssert = CSRFile_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_mstatus_prv = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  reg_mstatus_tsr = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  reg_mstatus_tw = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  reg_mstatus_tvm = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  reg_mstatus_mxr = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  reg_mstatus_sum = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  reg_mstatus_mprv = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  reg_mstatus_fs = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  reg_mstatus_mpp = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  reg_mstatus_spp = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  reg_mstatus_mpie = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  reg_mstatus_spie = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  reg_mstatus_mie = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  reg_mstatus_sie = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  reg_dcsr_prv = _RAND_14[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  reg_singleStepped = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  reg_dcsr_ebreakm = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  reg_dcsr_ebreaks = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  reg_dcsr_ebreaku = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  reg_debug = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{`RANDOM}};
  reg_mideleg = _RAND_20[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{`RANDOM}};
  reg_medeleg = _RAND_21[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  reg_dcsr_cause = _RAND_22[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  reg_dcsr_step = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {2{`RANDOM}};
  reg_dpc = _RAND_24[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {2{`RANDOM}};
  reg_dscratch = _RAND_25[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  reg_bp_0_control_dmode = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  reg_bp_0_control_action = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  reg_bp_0_control_tmatch = _RAND_28[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  reg_bp_0_control_m = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  reg_bp_0_control_s = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  reg_bp_0_control_u = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  reg_bp_0_control_x = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  reg_bp_0_control_w = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  reg_bp_0_control_r = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {2{`RANDOM}};
  reg_bp_0_address = _RAND_35[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  reg_pmp_0_cfg_l = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  reg_pmp_0_cfg_a = _RAND_37[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  reg_pmp_0_cfg_x = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  reg_pmp_0_cfg_w = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  reg_pmp_0_cfg_r = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  reg_pmp_0_addr = _RAND_41[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  reg_pmp_1_cfg_l = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  reg_pmp_1_cfg_a = _RAND_43[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  reg_pmp_1_cfg_x = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  reg_pmp_1_cfg_w = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  reg_pmp_1_cfg_r = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  reg_pmp_1_addr = _RAND_47[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  reg_pmp_2_cfg_l = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  reg_pmp_2_cfg_a = _RAND_49[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  reg_pmp_2_cfg_x = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  reg_pmp_2_cfg_w = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  reg_pmp_2_cfg_r = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  reg_pmp_2_addr = _RAND_53[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  reg_pmp_3_cfg_l = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  reg_pmp_3_cfg_a = _RAND_55[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  reg_pmp_3_cfg_x = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  reg_pmp_3_cfg_w = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  reg_pmp_3_cfg_r = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  reg_pmp_3_addr = _RAND_59[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  reg_pmp_4_cfg_l = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  reg_pmp_4_cfg_a = _RAND_61[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  reg_pmp_4_cfg_x = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  reg_pmp_4_cfg_w = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  reg_pmp_4_cfg_r = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  reg_pmp_4_addr = _RAND_65[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  reg_pmp_5_cfg_l = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  reg_pmp_5_cfg_a = _RAND_67[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  reg_pmp_5_cfg_x = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  reg_pmp_5_cfg_w = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  reg_pmp_5_cfg_r = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  reg_pmp_5_addr = _RAND_71[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  reg_pmp_6_cfg_l = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  reg_pmp_6_cfg_a = _RAND_73[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  reg_pmp_6_cfg_x = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  reg_pmp_6_cfg_w = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  reg_pmp_6_cfg_r = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  reg_pmp_6_addr = _RAND_77[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  reg_pmp_7_cfg_l = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  reg_pmp_7_cfg_a = _RAND_79[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  reg_pmp_7_cfg_x = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  reg_pmp_7_cfg_w = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  reg_pmp_7_cfg_r = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  reg_pmp_7_addr = _RAND_83[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {2{`RANDOM}};
  reg_mie = _RAND_84[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  reg_mip_seip = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  reg_mip_stip = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  reg_mip_ssip = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {2{`RANDOM}};
  reg_mepc = _RAND_88[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {2{`RANDOM}};
  reg_mcause = _RAND_89[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {2{`RANDOM}};
  reg_mbadaddr = _RAND_90[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {2{`RANDOM}};
  reg_mscratch = _RAND_91[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  reg_mtvec = _RAND_92[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  reg_mcounteren = _RAND_93[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  reg_scounteren = _RAND_94[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {2{`RANDOM}};
  reg_sepc = _RAND_95[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {2{`RANDOM}};
  reg_scause = _RAND_96[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {2{`RANDOM}};
  reg_sbadaddr = _RAND_97[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {2{`RANDOM}};
  reg_sscratch = _RAND_98[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {2{`RANDOM}};
  reg_stvec = _RAND_99[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  reg_sptbr_mode = _RAND_100[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {2{`RANDOM}};
  reg_sptbr_ppn = _RAND_101[43:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  reg_wfi = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  reg_fflags = _RAND_103[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  reg_frm = _RAND_104[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_286 = _RAND_105[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {2{`RANDOM}};
  _T_289 = _RAND_106[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_296 = _RAND_107[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {2{`RANDOM}};
  _T_299 = _RAND_108[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_310 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {2{`RANDOM}};
  reg_misa = _RAND_110[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  vpoffset_reg = _RAND_111[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  pcode_regs_0_locked = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  pcode_regs_1_locked = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  pcode_regs_2_locked = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  pcode_regs_3_locked = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  pcode_update_valid = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  pcode_update_bits_id = _RAND_117[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  pcode_update_bits_value_base = _RAND_118[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  pcode_update_bits_value_mask = _RAND_119[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  pcode_update_bits_value_valid = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  pcode_update_bits_value_locked = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  vpoffset_update_bits_value = _RAND_122[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_1626 = _RAND_123[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  CSRFile_state = _RAND_124[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    CSRFile_cov[initvar] = _RAND_125[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  CSRFile_covSum = _RAND_126[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  CSRFile_metaAssert = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      reg_mstatus_prv <= 2'h0;
    end else if (reset) begin
      reg_mstatus_prv <= 2'h3;
    end else if (_T_172) begin
      reg_mstatus_prv <= 2'h0;
    end else if (insn_ret) begin
      if (~io_rw_addr[9]) begin
        reg_mstatus_prv <= {{1'd0}, reg_mstatus_spp};
      end else if (io_rw_addr[10]) begin
        reg_mstatus_prv <= reg_dcsr_prv;
      end else begin
        reg_mstatus_prv <= reg_mstatus_mpp;
      end
    end else if (exception) begin
      if (trapToDebug) begin
        if (~reg_debug) begin
          reg_mstatus_prv <= 2'h3;
        end
      end else if (delegate) begin
        reg_mstatus_prv <= 2'h1;
      end else begin
        reg_mstatus_prv <= 2'h3;
      end
    end
    if (metaReset) begin
      reg_mstatus_tsr <= 1'h0;
    end else if (reset) begin
      reg_mstatus_tsr <= 1'h0;
    end else if (csr_wen) begin
      if (_T_983) begin
        reg_mstatus_tsr <= _T_3676[22];
      end
    end
    if (metaReset) begin
      reg_mstatus_tw <= 1'h0;
    end else if (reset) begin
      reg_mstatus_tw <= 1'h0;
    end else if (csr_wen) begin
      if (_T_983) begin
        reg_mstatus_tw <= _T_3676[21];
      end
    end
    if (metaReset) begin
      reg_mstatus_tvm <= 1'h0;
    end else if (reset) begin
      reg_mstatus_tvm <= 1'h0;
    end else if (csr_wen) begin
      if (_T_983) begin
        reg_mstatus_tvm <= _T_3676[20];
      end
    end
    if (metaReset) begin
      reg_mstatus_mxr <= 1'h0;
    end else if (reset) begin
      reg_mstatus_mxr <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1095) begin
        reg_mstatus_mxr <= _T_3676[19];
      end else if (_T_983) begin
        reg_mstatus_mxr <= _T_3676[19];
      end
    end
    if (metaReset) begin
      reg_mstatus_sum <= 1'h0;
    end else if (reset) begin
      reg_mstatus_sum <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1095) begin
        reg_mstatus_sum <= _T_3676[18];
      end else if (_T_983) begin
        reg_mstatus_sum <= _T_3676[18];
      end
    end
    if (metaReset) begin
      reg_mstatus_mprv <= 1'h0;
    end else if (reset) begin
      reg_mstatus_mprv <= 1'h0;
    end else if (csr_wen) begin
      if (_T_983) begin
        reg_mstatus_mprv <= _T_3676[17];
      end
    end
    if (metaReset) begin
      reg_mstatus_fs <= 2'h0;
    end else if (reset) begin
      reg_mstatus_fs <= 2'h0;
    end else if (csr_wen) begin
      if (_T_1095) begin
        if (_T_3708) begin
          reg_mstatus_fs <= 2'h3;
        end else begin
          reg_mstatus_fs <= 2'h0;
        end
      end else if (_T_983) begin
        if (_T_3708) begin
          reg_mstatus_fs <= 2'h3;
        end else begin
          reg_mstatus_fs <= 2'h0;
        end
      end
    end
    if (metaReset) begin
      reg_mstatus_mpp <= 2'h0;
    end else if (reset) begin
      reg_mstatus_mpp <= 2'h3;
    end else if (csr_wen) begin
      if (_T_983) begin
        if (_T_3706) begin
          reg_mstatus_mpp <= 2'h0;
        end else begin
          reg_mstatus_mpp <= _T_3676[12:11];
        end
      end else if (insn_ret) begin
        if (~io_rw_addr[9]) begin
          if (exception) begin
            if (!(trapToDebug)) begin
              if (!(delegate)) begin
                reg_mstatus_mpp <= reg_mstatus_prv;
              end
            end
          end
        end else if (io_rw_addr[10]) begin
          if (exception) begin
            if (!(trapToDebug)) begin
              if (!(delegate)) begin
                reg_mstatus_mpp <= reg_mstatus_prv;
              end
            end
          end
        end else begin
          reg_mstatus_mpp <= 2'h0;
        end
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (!(delegate)) begin
            reg_mstatus_mpp <= reg_mstatus_prv;
          end
        end
      end
    end else if (insn_ret) begin
      if (~io_rw_addr[9]) begin
        if (exception) begin
          if (!(trapToDebug)) begin
            if (!(delegate)) begin
              reg_mstatus_mpp <= reg_mstatus_prv;
            end
          end
        end
      end else if (io_rw_addr[10]) begin
        reg_mstatus_mpp <= _GEN_123;
      end else begin
        reg_mstatus_mpp <= 2'h0;
      end
    end else begin
      reg_mstatus_mpp <= _GEN_123;
    end
    if (metaReset) begin
      reg_mstatus_spp <= 1'h0;
    end else if (reset) begin
      reg_mstatus_spp <= 1'h0;
    end else begin
      reg_mstatus_spp <= _GEN_562[0];
    end
    if (metaReset) begin
      reg_mstatus_mpie <= 1'h0;
    end else if (reset) begin
      reg_mstatus_mpie <= 1'h0;
    end else if (csr_wen) begin
      if (_T_983) begin
        reg_mstatus_mpie <= _T_3676[7];
      end else if (insn_ret) begin
        if (~io_rw_addr[9]) begin
          if (exception) begin
            if (!(trapToDebug)) begin
              if (!(delegate)) begin
                reg_mstatus_mpie <= reg_mstatus_mie;
              end
            end
          end
        end else if (io_rw_addr[10]) begin
          if (exception) begin
            if (!(trapToDebug)) begin
              if (!(delegate)) begin
                reg_mstatus_mpie <= reg_mstatus_mie;
              end
            end
          end
        end else begin
          reg_mstatus_mpie <= 1'h1;
        end
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (!(delegate)) begin
            reg_mstatus_mpie <= reg_mstatus_mie;
          end
        end
      end
    end else if (insn_ret) begin
      if (~io_rw_addr[9]) begin
        if (exception) begin
          if (!(trapToDebug)) begin
            if (!(delegate)) begin
              reg_mstatus_mpie <= reg_mstatus_mie;
            end
          end
        end
      end else if (io_rw_addr[10]) begin
        reg_mstatus_mpie <= _GEN_122;
      end else begin
        reg_mstatus_mpie <= 1'h1;
      end
    end else begin
      reg_mstatus_mpie <= _GEN_122;
    end
    if (metaReset) begin
      reg_mstatus_spie <= 1'h0;
    end else if (reset) begin
      reg_mstatus_spie <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1095) begin
        reg_mstatus_spie <= _T_3676[5];
      end else if (_T_983) begin
        reg_mstatus_spie <= _T_3676[5];
      end else if (insn_ret) begin
        reg_mstatus_spie <= _GEN_132;
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (delegate) begin
            reg_mstatus_spie <= reg_mstatus_sie;
          end
        end
      end
    end else if (insn_ret) begin
      reg_mstatus_spie <= _GEN_132;
    end else if (exception) begin
      if (!(trapToDebug)) begin
        if (delegate) begin
          reg_mstatus_spie <= reg_mstatus_sie;
        end
      end
    end
    if (metaReset) begin
      reg_mstatus_mie <= 1'h0;
    end else if (reset) begin
      reg_mstatus_mie <= 1'h0;
    end else if (csr_wen) begin
      if (_T_983) begin
        reg_mstatus_mie <= _T_3676[3];
      end else if (insn_ret) begin
        if (~io_rw_addr[9]) begin
          if (exception) begin
            if (!(trapToDebug)) begin
              reg_mstatus_mie <= _GEN_88;
            end
          end
        end else if (io_rw_addr[10]) begin
          if (exception) begin
            if (!(trapToDebug)) begin
              reg_mstatus_mie <= _GEN_88;
            end
          end
        end else begin
          reg_mstatus_mie <= reg_mstatus_mpie;
        end
      end else if (exception) begin
        if (!(trapToDebug)) begin
          reg_mstatus_mie <= _GEN_88;
        end
      end
    end else if (insn_ret) begin
      if (~io_rw_addr[9]) begin
        if (exception) begin
          if (!(trapToDebug)) begin
            reg_mstatus_mie <= _GEN_88;
          end
        end
      end else if (io_rw_addr[10]) begin
        reg_mstatus_mie <= _GEN_124;
      end else begin
        reg_mstatus_mie <= reg_mstatus_mpie;
      end
    end else begin
      reg_mstatus_mie <= _GEN_124;
    end
    if (metaReset) begin
      reg_mstatus_sie <= 1'h0;
    end else if (reset) begin
      reg_mstatus_sie <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1095) begin
        reg_mstatus_sie <= _T_3676[1];
      end else if (_T_983) begin
        reg_mstatus_sie <= _T_3676[1];
      end else if (insn_ret) begin
        if (~io_rw_addr[9]) begin
          reg_mstatus_sie <= reg_mstatus_spie;
        end else if (exception) begin
          if (!(trapToDebug)) begin
            if (delegate) begin
              reg_mstatus_sie <= 1'h0;
            end
          end
        end
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (delegate) begin
            reg_mstatus_sie <= 1'h0;
          end
        end
      end
    end else if (insn_ret) begin
      if (~io_rw_addr[9]) begin
        reg_mstatus_sie <= reg_mstatus_spie;
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (delegate) begin
            reg_mstatus_sie <= 1'h0;
          end
        end
      end
    end else if (exception) begin
      if (!(trapToDebug)) begin
        if (delegate) begin
          reg_mstatus_sie <= 1'h0;
        end
      end
    end
    if (metaReset) begin
      reg_dcsr_prv <= 2'h0;
    end else if (reset) begin
      reg_dcsr_prv <= 2'h3;
    end else if (csr_wen) begin
      if (_T_992) begin
        if (_T_3813) begin
          reg_dcsr_prv <= 2'h0;
        end else begin
          reg_dcsr_prv <= wdata[1:0];
        end
      end else if (exception) begin
        if (trapToDebug) begin
          if (~reg_debug) begin
            reg_dcsr_prv <= reg_mstatus_prv;
          end
        end
      end
    end else if (exception) begin
      if (trapToDebug) begin
        if (~reg_debug) begin
          reg_dcsr_prv <= reg_mstatus_prv;
        end
      end
    end
    if (metaReset) begin
      reg_singleStepped <= 1'h0;
    end else if (~io_singleStep) begin
      reg_singleStepped <= 1'h0;
    end else begin
      reg_singleStepped <= _GEN_68;
    end
    if (metaReset) begin
      reg_dcsr_ebreakm <= 1'h0;
    end else if (reset) begin
      reg_dcsr_ebreakm <= 1'h0;
    end else if (csr_wen) begin
      if (_T_992) begin
        reg_dcsr_ebreakm <= wdata[15];
      end
    end
    if (metaReset) begin
      reg_dcsr_ebreaks <= 1'h0;
    end else if (reset) begin
      reg_dcsr_ebreaks <= 1'h0;
    end else if (csr_wen) begin
      if (_T_992) begin
        reg_dcsr_ebreaks <= wdata[13];
      end
    end
    if (metaReset) begin
      reg_dcsr_ebreaku <= 1'h0;
    end else if (reset) begin
      reg_dcsr_ebreaku <= 1'h0;
    end else if (csr_wen) begin
      if (_T_992) begin
        reg_dcsr_ebreaku <= wdata[12];
      end
    end
    if (metaReset) begin
      reg_debug <= 1'h0;
    end else if (reset) begin
      reg_debug <= 1'h0;
    end else if (insn_ret) begin
      if (~io_rw_addr[9]) begin
        if (exception) begin
          if (trapToDebug) begin
            reg_debug <= _GEN_70;
          end
        end
      end else if (io_rw_addr[10]) begin
        reg_debug <= 1'h0;
      end else if (exception) begin
        if (trapToDebug) begin
          reg_debug <= _GEN_70;
        end
      end
    end else if (exception) begin
      if (trapToDebug) begin
        reg_debug <= _GEN_70;
      end
    end
    if (metaReset) begin
      reg_mideleg <= 64'h0;
    end else if (csr_wen) begin
      if (_T_1105) begin
        reg_mideleg <= _T_3915;
      end
    end
    if (metaReset) begin
      reg_medeleg <= 64'h0;
    end else if (csr_wen) begin
      if (_T_1106) begin
        reg_medeleg <= _T_3916;
      end
    end
    if (metaReset) begin
      reg_dcsr_cause <= 3'h0;
    end else if (reset) begin
      reg_dcsr_cause <= 3'h0;
    end else if (exception) begin
      if (trapToDebug) begin
        if (~reg_debug) begin
          if (reg_singleStepped) begin
            reg_dcsr_cause <= 3'h4;
          end else begin
            reg_dcsr_cause <= {{1'd0}, _T_1662};
          end
        end
      end
    end
    if (metaReset) begin
      reg_dcsr_step <= 1'h0;
    end else if (reset) begin
      reg_dcsr_step <= 1'h0;
    end else if (csr_wen) begin
      if (_T_992) begin
        reg_dcsr_step <= wdata[2];
      end
    end
    if (metaReset) begin
      reg_dpc <= 40'h0;
    end else begin
      reg_dpc <= _GEN_591[39:0];
    end
    if (metaReset) begin
      reg_dscratch <= 64'h0;
    end else if (csr_wen) begin
      if (_T_994) begin
        reg_dscratch <= wdata;
      end
    end
    if (metaReset) begin
      reg_bp_0_control_dmode <= 1'h0;
    end else if (reset) begin
      reg_bp_0_control_dmode <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3921) begin
        if (_T_980) begin
          reg_bp_0_control_dmode <= _T_3942;
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_action <= 1'h0;
    end else if (reset) begin
      reg_bp_0_control_action <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3921) begin
        if (_T_980) begin
          reg_bp_0_control_action <= _T_3943;
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_tmatch <= 2'h0;
    end else if (csr_wen) begin
      if (_T_3921) begin
        if (_T_980) begin
          reg_bp_0_control_tmatch <= wdata[8:7];
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_m <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3921) begin
        if (_T_980) begin
          reg_bp_0_control_m <= wdata[6];
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_s <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3921) begin
        if (_T_980) begin
          reg_bp_0_control_s <= wdata[4];
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_u <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3921) begin
        if (_T_980) begin
          reg_bp_0_control_u <= wdata[3];
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_x <= 1'h0;
    end else if (reset) begin
      reg_bp_0_control_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3921) begin
        if (_T_980) begin
          reg_bp_0_control_x <= wdata[2];
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_w <= 1'h0;
    end else if (reset) begin
      reg_bp_0_control_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3921) begin
        if (_T_980) begin
          reg_bp_0_control_w <= wdata[1];
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_r <= 1'h0;
    end else if (reset) begin
      reg_bp_0_control_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3921) begin
        if (_T_980) begin
          reg_bp_0_control_r <= wdata[0];
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_address <= 39'h0;
    end else if (csr_wen) begin
      if (_T_3921) begin
        if (_T_981) begin
          reg_bp_0_address <= wdata[38:0];
        end
      end
    end
    if (metaReset) begin
      reg_pmp_0_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_0_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3945) begin
        reg_pmp_0_cfg_l <= wdata[7];
      end
    end
    if (metaReset) begin
      reg_pmp_0_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_0_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_3945) begin
        reg_pmp_0_cfg_a <= wdata[4:3];
      end
    end
    if (metaReset) begin
      reg_pmp_0_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3945) begin
        reg_pmp_0_cfg_x <= wdata[2];
      end
    end
    if (metaReset) begin
      reg_pmp_0_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3945) begin
        reg_pmp_0_cfg_w <= wdata[1];
      end
    end
    if (metaReset) begin
      reg_pmp_0_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3945) begin
        reg_pmp_0_cfg_r <= wdata[0];
      end
    end
    if (metaReset) begin
      reg_pmp_0_addr <= 30'h0;
    end else begin
      reg_pmp_0_addr <= _GEN_643[29:0];
    end
    if (metaReset) begin
      reg_pmp_1_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_1_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3967) begin
        reg_pmp_1_cfg_l <= wdata[15];
      end
    end
    if (metaReset) begin
      reg_pmp_1_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_1_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_3967) begin
        reg_pmp_1_cfg_a <= wdata[12:11];
      end
    end
    if (metaReset) begin
      reg_pmp_1_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3967) begin
        reg_pmp_1_cfg_x <= wdata[10];
      end
    end
    if (metaReset) begin
      reg_pmp_1_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3967) begin
        reg_pmp_1_cfg_w <= wdata[9];
      end
    end
    if (metaReset) begin
      reg_pmp_1_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3967) begin
        reg_pmp_1_cfg_r <= wdata[8];
      end
    end
    if (metaReset) begin
      reg_pmp_1_addr <= 30'h0;
    end else begin
      reg_pmp_1_addr <= _GEN_650[29:0];
    end
    if (metaReset) begin
      reg_pmp_2_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_2_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3989) begin
        reg_pmp_2_cfg_l <= wdata[23];
      end
    end
    if (metaReset) begin
      reg_pmp_2_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_2_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_3989) begin
        reg_pmp_2_cfg_a <= wdata[20:19];
      end
    end
    if (metaReset) begin
      reg_pmp_2_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3989) begin
        reg_pmp_2_cfg_x <= wdata[18];
      end
    end
    if (metaReset) begin
      reg_pmp_2_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3989) begin
        reg_pmp_2_cfg_w <= wdata[17];
      end
    end
    if (metaReset) begin
      reg_pmp_2_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_3989) begin
        reg_pmp_2_cfg_r <= wdata[16];
      end
    end
    if (metaReset) begin
      reg_pmp_2_addr <= 30'h0;
    end else begin
      reg_pmp_2_addr <= _GEN_657[29:0];
    end
    if (metaReset) begin
      reg_pmp_3_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_3_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4011) begin
        reg_pmp_3_cfg_l <= wdata[31];
      end
    end
    if (metaReset) begin
      reg_pmp_3_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_3_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_4011) begin
        reg_pmp_3_cfg_a <= wdata[28:27];
      end
    end
    if (metaReset) begin
      reg_pmp_3_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4011) begin
        reg_pmp_3_cfg_x <= wdata[26];
      end
    end
    if (metaReset) begin
      reg_pmp_3_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4011) begin
        reg_pmp_3_cfg_w <= wdata[25];
      end
    end
    if (metaReset) begin
      reg_pmp_3_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4011) begin
        reg_pmp_3_cfg_r <= wdata[24];
      end
    end
    if (metaReset) begin
      reg_pmp_3_addr <= 30'h0;
    end else begin
      reg_pmp_3_addr <= _GEN_664[29:0];
    end
    if (metaReset) begin
      reg_pmp_4_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_4_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4033) begin
        reg_pmp_4_cfg_l <= wdata[39];
      end
    end
    if (metaReset) begin
      reg_pmp_4_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_4_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_4033) begin
        reg_pmp_4_cfg_a <= wdata[36:35];
      end
    end
    if (metaReset) begin
      reg_pmp_4_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4033) begin
        reg_pmp_4_cfg_x <= wdata[34];
      end
    end
    if (metaReset) begin
      reg_pmp_4_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4033) begin
        reg_pmp_4_cfg_w <= wdata[33];
      end
    end
    if (metaReset) begin
      reg_pmp_4_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4033) begin
        reg_pmp_4_cfg_r <= wdata[32];
      end
    end
    if (metaReset) begin
      reg_pmp_4_addr <= 30'h0;
    end else begin
      reg_pmp_4_addr <= _GEN_671[29:0];
    end
    if (metaReset) begin
      reg_pmp_5_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_5_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4055) begin
        reg_pmp_5_cfg_l <= wdata[47];
      end
    end
    if (metaReset) begin
      reg_pmp_5_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_5_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_4055) begin
        reg_pmp_5_cfg_a <= wdata[44:43];
      end
    end
    if (metaReset) begin
      reg_pmp_5_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4055) begin
        reg_pmp_5_cfg_x <= wdata[42];
      end
    end
    if (metaReset) begin
      reg_pmp_5_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4055) begin
        reg_pmp_5_cfg_w <= wdata[41];
      end
    end
    if (metaReset) begin
      reg_pmp_5_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4055) begin
        reg_pmp_5_cfg_r <= wdata[40];
      end
    end
    if (metaReset) begin
      reg_pmp_5_addr <= 30'h0;
    end else begin
      reg_pmp_5_addr <= _GEN_678[29:0];
    end
    if (metaReset) begin
      reg_pmp_6_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_6_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4077) begin
        reg_pmp_6_cfg_l <= wdata[55];
      end
    end
    if (metaReset) begin
      reg_pmp_6_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_6_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_4077) begin
        reg_pmp_6_cfg_a <= wdata[52:51];
      end
    end
    if (metaReset) begin
      reg_pmp_6_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4077) begin
        reg_pmp_6_cfg_x <= wdata[50];
      end
    end
    if (metaReset) begin
      reg_pmp_6_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4077) begin
        reg_pmp_6_cfg_w <= wdata[49];
      end
    end
    if (metaReset) begin
      reg_pmp_6_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4077) begin
        reg_pmp_6_cfg_r <= wdata[48];
      end
    end
    if (metaReset) begin
      reg_pmp_6_addr <= 30'h0;
    end else begin
      reg_pmp_6_addr <= _GEN_685[29:0];
    end
    if (metaReset) begin
      reg_pmp_7_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_7_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4099) begin
        reg_pmp_7_cfg_l <= wdata[63];
      end
    end
    if (metaReset) begin
      reg_pmp_7_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_7_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_4099) begin
        reg_pmp_7_cfg_a <= wdata[60:59];
      end
    end
    if (metaReset) begin
      reg_pmp_7_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4099) begin
        reg_pmp_7_cfg_x <= wdata[58];
      end
    end
    if (metaReset) begin
      reg_pmp_7_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4099) begin
        reg_pmp_7_cfg_w <= wdata[57];
      end
    end
    if (metaReset) begin
      reg_pmp_7_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_4099) begin
        reg_pmp_7_cfg_r <= wdata[56];
      end
    end
    if (metaReset) begin
      reg_pmp_7_addr <= 30'h0;
    end else begin
      reg_pmp_7_addr <= _GEN_692[29:0];
    end
    if (metaReset) begin
      reg_mie <= 64'h0;
    end else if (csr_wen) begin
      if (_T_1097) begin
        reg_mie <= _T_3903;
      end else if (_T_986) begin
        reg_mie <= _T_3777;
      end
    end
    if (metaReset) begin
      reg_mip_seip <= 1'h0;
    end else if (csr_wen) begin
      if (_T_985) begin
        reg_mip_seip <= _T_3749[9];
      end
    end
    if (metaReset) begin
      reg_mip_stip <= 1'h0;
    end else if (csr_wen) begin
      if (_T_985) begin
        reg_mip_stip <= _T_3749[5];
      end
    end
    if (metaReset) begin
      reg_mip_ssip <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1096) begin
        reg_mip_ssip <= _T_3861[1];
      end else if (_T_985) begin
        reg_mip_ssip <= _T_3749[1];
      end
    end
    if (metaReset) begin
      reg_mepc <= 40'h0;
    end else begin
      reg_mepc <= _GEN_574[39:0];
    end
    if (metaReset) begin
      reg_mcause <= 64'h0;
    end else if (csr_wen) begin
      if (_T_990) begin
        reg_mcause <= _T_3787;
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (!(delegate)) begin
            if (insn_call) begin
              reg_mcause <= {{60'd0}, _T_1572};
            end else if (insn_break) begin
              reg_mcause <= 64'h3;
            end else begin
              reg_mcause <= io_cause;
            end
          end
        end
      end
    end else if (exception) begin
      if (!(trapToDebug)) begin
        if (!(delegate)) begin
          if (insn_call) begin
            reg_mcause <= {{60'd0}, _T_1572};
          end else if (insn_break) begin
            reg_mcause <= 64'h3;
          end else begin
            reg_mcause <= io_cause;
          end
        end
      end
    end
    if (metaReset) begin
      reg_mbadaddr <= 40'h0;
    end else if (csr_wen) begin
      if (_T_989) begin
        reg_mbadaddr <= wdata[39:0];
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (!(delegate)) begin
            reg_mbadaddr <= io_tval;
          end
        end
      end
    end else if (exception) begin
      if (!(trapToDebug)) begin
        if (!(delegate)) begin
          reg_mbadaddr <= io_tval;
        end
      end
    end
    if (metaReset) begin
      reg_mscratch <= 64'h0;
    end else if (csr_wen) begin
      if (_T_987) begin
        reg_mscratch <= wdata;
      end
    end
    if (metaReset) begin
      reg_mtvec <= 32'h0;
    end else if (reset) begin
      reg_mtvec <= 32'h0;
    end else begin
      reg_mtvec <= _GEN_576[31:0];
    end
    if (metaReset) begin
      reg_mcounteren <= 32'h0;
    end else begin
      reg_mcounteren <= _GEN_603[31:0];
    end
    if (metaReset) begin
      reg_scounteren <= 32'h0;
    end else begin
      reg_scounteren <= _GEN_602[31:0];
    end
    if (metaReset) begin
      reg_sepc <= 40'h0;
    end else begin
      reg_sepc <= _GEN_596[39:0];
    end
    if (metaReset) begin
      reg_scause <= 64'h0;
    end else if (csr_wen) begin
      if (_T_1099) begin
        reg_scause <= _T_3913;
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (delegate) begin
            if (insn_call) begin
              reg_scause <= {{60'd0}, _T_1572};
            end else if (insn_break) begin
              reg_scause <= 64'h3;
            end else begin
              reg_scause <= io_cause;
            end
          end
        end
      end
    end else if (exception) begin
      if (!(trapToDebug)) begin
        if (delegate) begin
          if (insn_call) begin
            reg_scause <= {{60'd0}, _T_1572};
          end else if (insn_break) begin
            reg_scause <= 64'h3;
          end else begin
            reg_scause <= io_cause;
          end
        end
      end
    end
    if (metaReset) begin
      reg_sbadaddr <= 40'h0;
    end else if (csr_wen) begin
      if (_T_1100) begin
        reg_sbadaddr <= wdata[39:0];
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (delegate) begin
            reg_sbadaddr <= io_tval;
          end
        end
      end
    end else if (exception) begin
      if (!(trapToDebug)) begin
        if (delegate) begin
          reg_sbadaddr <= io_tval;
        end
      end
    end
    if (metaReset) begin
      reg_sscratch <= 64'h0;
    end else if (csr_wen) begin
      if (_T_1098) begin
        reg_sscratch <= wdata;
      end
    end
    if (metaReset) begin
      reg_stvec <= 39'h0;
    end else begin
      reg_stvec <= _GEN_597[38:0];
    end
    if (metaReset) begin
      reg_sptbr_mode <= 4'h0;
    end else if (csr_wen) begin
      if (_T_1101) begin
        if (_T_3895) begin
          reg_sptbr_mode <= 4'h8;
        end else if (_T_3894) begin
          reg_sptbr_mode <= 4'h0;
        end
      end
    end
    if (metaReset) begin
      reg_sptbr_ppn <= 44'h0;
    end else if (csr_wen) begin
      if (_T_1101) begin
        if (_T_3898) begin
          reg_sptbr_ppn <= {{24'd0}, wdata[19:0]};
        end
      end
    end
    if (metaReset) begin
      reg_fflags <= 5'h0;
    end else begin
      reg_fflags <= _GEN_584[4:0];
    end
    if (metaReset) begin
      reg_frm <= 3'h0;
    end else begin
      reg_frm <= _GEN_585[2:0];
    end
    if (metaReset) begin
      _T_286 <= 6'h0;
    end else if (reset) begin
      _T_286 <= 6'h0;
    end else begin
      _T_286 <= _GEN_581[5:0];
    end
    if (metaReset) begin
      _T_289 <= 58'h0;
    end else if (reset) begin
      _T_289 <= 58'h0;
    end else if (csr_wen) begin
      if (_T_999) begin
        _T_289 <= wdata[63:6];
      end else if (_T_287[6]) begin
        _T_289 <= _T_292;
      end
    end else if (_T_287[6]) begin
      _T_289 <= _T_292;
    end
    if (metaReset) begin
      _T_310 <= 1'h0;
    end else begin
      _T_310 <= io_interrupts_seip;
    end
    if (metaReset) begin
      reg_misa <= 64'h0;
    end else if (reset) begin
      reg_misa <= 64'h800000000014112d;
    end else if (csr_wen) begin
      if (_T_982) begin
        if (_T_3716) begin
          reg_misa <= _T_3725;
        end
      end
    end
    if (metaReset) begin
      vpoffset_reg <= 27'h0;
    end else if (csr_wen) begin
      if (_T_1090) begin
        vpoffset_reg <= wdata[38:12];
      end
    end
    if (metaReset) begin
      pcode_regs_0_locked <= 1'h0;
    end else if (reset) begin
      pcode_regs_0_locked <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1091) begin
        if (~pcode_regs_0_locked) begin
          pcode_regs_0_locked <= wdata[0];
        end
      end
    end
    if (metaReset) begin
      pcode_regs_1_locked <= 1'h0;
    end else if (reset) begin
      pcode_regs_1_locked <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1092) begin
        if (~pcode_regs_1_locked) begin
          pcode_regs_1_locked <= wdata[0];
        end
      end
    end
    if (metaReset) begin
      pcode_regs_2_locked <= 1'h0;
    end else if (reset) begin
      pcode_regs_2_locked <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1093) begin
        if (~pcode_regs_2_locked) begin
          pcode_regs_2_locked <= wdata[0];
        end
      end
    end
    if (metaReset) begin
      pcode_regs_3_locked <= 1'h0;
    end else if (reset) begin
      pcode_regs_3_locked <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1094) begin
        if (~pcode_regs_3_locked) begin
          pcode_regs_3_locked <= wdata[0];
        end
      end
    end
    if (metaReset) begin
      pcode_update_valid <= 1'h0;
    end else begin
      pcode_update_valid <= csr_wen & _GEN_304;
    end
    if (metaReset) begin
      pcode_update_bits_id <= 2'h0;
    end else begin
      pcode_update_bits_id <= _GEN_547[1:0];
    end
    if (metaReset) begin
      pcode_update_bits_value_base <= 20'h0;
    end else if (csr_wen) begin
      if (_T_1094) begin
        if (~pcode_regs_3_locked) begin
          pcode_update_bits_value_base <= wdata[31:12];
        end else if (_T_1093) begin
          if (~pcode_regs_2_locked) begin
            pcode_update_bits_value_base <= wdata[31:12];
          end else if (_T_1092) begin
            if (~pcode_regs_1_locked) begin
              pcode_update_bits_value_base <= wdata[31:12];
            end else if (_T_1091) begin
              if (~pcode_regs_0_locked) begin
                pcode_update_bits_value_base <= wdata[31:12];
              end
            end
          end else if (_T_1091) begin
            if (~pcode_regs_0_locked) begin
              pcode_update_bits_value_base <= wdata[31:12];
            end
          end
        end else if (_T_1092) begin
          if (~pcode_regs_1_locked) begin
            pcode_update_bits_value_base <= wdata[31:12];
          end else if (_T_1091) begin
            if (~pcode_regs_0_locked) begin
              pcode_update_bits_value_base <= wdata[31:12];
            end
          end
        end else if (_T_1091) begin
          if (~pcode_regs_0_locked) begin
            pcode_update_bits_value_base <= wdata[31:12];
          end
        end
      end else if (_T_1093) begin
        if (~pcode_regs_2_locked) begin
          pcode_update_bits_value_base <= wdata[31:12];
        end else if (_T_1092) begin
          if (~pcode_regs_1_locked) begin
            pcode_update_bits_value_base <= wdata[31:12];
          end else begin
            pcode_update_bits_value_base <= _GEN_186;
          end
        end else begin
          pcode_update_bits_value_base <= _GEN_186;
        end
      end else if (_T_1092) begin
        if (~pcode_regs_1_locked) begin
          pcode_update_bits_value_base <= wdata[31:12];
        end else begin
          pcode_update_bits_value_base <= _GEN_186;
        end
      end else begin
        pcode_update_bits_value_base <= _GEN_186;
      end
    end
    if (metaReset) begin
      pcode_update_bits_value_mask <= 10'h0;
    end else if (csr_wen) begin
      if (_T_1094) begin
        if (~pcode_regs_3_locked) begin
          pcode_update_bits_value_mask <= wdata[11:2];
        end else if (_T_1093) begin
          if (~pcode_regs_2_locked) begin
            pcode_update_bits_value_mask <= wdata[11:2];
          end else if (_T_1092) begin
            if (~pcode_regs_1_locked) begin
              pcode_update_bits_value_mask <= wdata[11:2];
            end else if (_T_1091) begin
              if (~pcode_regs_0_locked) begin
                pcode_update_bits_value_mask <= wdata[11:2];
              end
            end
          end else if (_T_1091) begin
            if (~pcode_regs_0_locked) begin
              pcode_update_bits_value_mask <= wdata[11:2];
            end
          end
        end else if (_T_1092) begin
          if (~pcode_regs_1_locked) begin
            pcode_update_bits_value_mask <= wdata[11:2];
          end else if (_T_1091) begin
            if (~pcode_regs_0_locked) begin
              pcode_update_bits_value_mask <= wdata[11:2];
            end
          end
        end else if (_T_1091) begin
          if (~pcode_regs_0_locked) begin
            pcode_update_bits_value_mask <= wdata[11:2];
          end
        end
      end else if (_T_1093) begin
        if (~pcode_regs_2_locked) begin
          pcode_update_bits_value_mask <= wdata[11:2];
        end else if (_T_1092) begin
          if (~pcode_regs_1_locked) begin
            pcode_update_bits_value_mask <= wdata[11:2];
          end else begin
            pcode_update_bits_value_mask <= _GEN_187;
          end
        end else begin
          pcode_update_bits_value_mask <= _GEN_187;
        end
      end else if (_T_1092) begin
        if (~pcode_regs_1_locked) begin
          pcode_update_bits_value_mask <= wdata[11:2];
        end else begin
          pcode_update_bits_value_mask <= _GEN_187;
        end
      end else begin
        pcode_update_bits_value_mask <= _GEN_187;
      end
    end
    if (metaReset) begin
      pcode_update_bits_value_valid <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1094) begin
        if (~pcode_regs_3_locked) begin
          pcode_update_bits_value_valid <= wdata[1];
        end else if (_T_1093) begin
          if (~pcode_regs_2_locked) begin
            pcode_update_bits_value_valid <= wdata[1];
          end else if (_T_1092) begin
            if (~pcode_regs_1_locked) begin
              pcode_update_bits_value_valid <= wdata[1];
            end else if (_T_1091) begin
              if (~pcode_regs_0_locked) begin
                pcode_update_bits_value_valid <= wdata[1];
              end
            end
          end else if (_T_1091) begin
            if (~pcode_regs_0_locked) begin
              pcode_update_bits_value_valid <= wdata[1];
            end
          end
        end else if (_T_1092) begin
          if (~pcode_regs_1_locked) begin
            pcode_update_bits_value_valid <= wdata[1];
          end else if (_T_1091) begin
            if (~pcode_regs_0_locked) begin
              pcode_update_bits_value_valid <= wdata[1];
            end
          end
        end else if (_T_1091) begin
          if (~pcode_regs_0_locked) begin
            pcode_update_bits_value_valid <= wdata[1];
          end
        end
      end else if (_T_1093) begin
        if (~pcode_regs_2_locked) begin
          pcode_update_bits_value_valid <= wdata[1];
        end else if (_T_1092) begin
          if (~pcode_regs_1_locked) begin
            pcode_update_bits_value_valid <= wdata[1];
          end else begin
            pcode_update_bits_value_valid <= _GEN_188;
          end
        end else begin
          pcode_update_bits_value_valid <= _GEN_188;
        end
      end else if (_T_1092) begin
        if (~pcode_regs_1_locked) begin
          pcode_update_bits_value_valid <= wdata[1];
        end else begin
          pcode_update_bits_value_valid <= _GEN_188;
        end
      end else begin
        pcode_update_bits_value_valid <= _GEN_188;
      end
    end
    if (metaReset) begin
      pcode_update_bits_value_locked <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1094) begin
        if (~pcode_regs_3_locked) begin
          pcode_update_bits_value_locked <= wdata[0];
        end else if (_T_1093) begin
          if (~pcode_regs_2_locked) begin
            pcode_update_bits_value_locked <= wdata[0];
          end else if (_T_1092) begin
            if (~pcode_regs_1_locked) begin
              pcode_update_bits_value_locked <= wdata[0];
            end else if (_T_1091) begin
              if (~pcode_regs_0_locked) begin
                pcode_update_bits_value_locked <= wdata[0];
              end
            end
          end else if (_T_1091) begin
            if (~pcode_regs_0_locked) begin
              pcode_update_bits_value_locked <= wdata[0];
            end
          end
        end else if (_T_1092) begin
          if (~pcode_regs_1_locked) begin
            pcode_update_bits_value_locked <= wdata[0];
          end else if (_T_1091) begin
            if (~pcode_regs_0_locked) begin
              pcode_update_bits_value_locked <= wdata[0];
            end
          end
        end else if (_T_1091) begin
          if (~pcode_regs_0_locked) begin
            pcode_update_bits_value_locked <= wdata[0];
          end
        end
      end else if (_T_1093) begin
        if (~pcode_regs_2_locked) begin
          pcode_update_bits_value_locked <= wdata[0];
        end else if (_T_1092) begin
          if (~pcode_regs_1_locked) begin
            pcode_update_bits_value_locked <= wdata[0];
          end else begin
            pcode_update_bits_value_locked <= _GEN_189;
          end
        end else begin
          pcode_update_bits_value_locked <= _GEN_189;
        end
      end else if (_T_1092) begin
        if (~pcode_regs_1_locked) begin
          pcode_update_bits_value_locked <= wdata[0];
        end else begin
          pcode_update_bits_value_locked <= _GEN_189;
        end
      end else begin
        pcode_update_bits_value_locked <= _GEN_189;
      end
    end
    if (metaReset) begin
      vpoffset_update_bits_value <= 27'h0;
    end else if (csr_wen) begin
      if (_T_1090) begin
        vpoffset_update_bits_value <= wdata[38:12];
      end
    end
    if (metaReset) begin
      _T_1626 <= 2'h0;
    end else if (_T_1623) begin
      _T_1626 <= reg_mstatus_mpp;
    end else begin
      _T_1626 <= reg_mstatus_prv;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_1633) begin
          $fwrite(32'h80000002,"Assertion failed: these conditions must be mutually exclusive\n    at CSR.scala:656 assert(PopCount(insn_ret :: insn_call :: insn_break :: io.exception :: Nil) <= 1, \"these conditions must be mutually exclusive\")\n"); // @[CSR.scala 656:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_1633) begin
          $fatal; // @[CSR.scala 656:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_1655) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CSR.scala:664 assert(!reg_singleStepped || io.retire === UInt(0))\n"); // @[CSR.scala 664:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_1655) begin
          $fatal; // @[CSR.scala 664:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    CSRFile_state <= CSRFile_xor0;
    if (!(CSRFile_cov_read_data)) begin
      CSRFile_covSum <= CSRFile_covSum + 1'h1;
    end
    if (metaReset) begin
      CSRFile_metaAssert <= 1'h0;
    end else begin
      CSRFile_metaAssert <= CSRFile_metaAssert | CSRFile_or0;
    end
  end
  always @(posedge io_ungated_clock) begin
    if (metaReset) begin
      reg_wfi <= 1'h0;
    end else if (reset) begin
      reg_wfi <= 1'h0;
    end else if (_T_1641) begin
      reg_wfi <= 1'h0;
    end else begin
      reg_wfi <= _GEN_66;
    end
    if (metaReset) begin
      _T_296 <= 6'h0;
    end else if (reset) begin
      _T_296 <= 6'h0;
    end else begin
      _T_296 <= _GEN_579[5:0];
    end
    if (metaReset) begin
      _T_299 <= 58'h0;
    end else if (reset) begin
      _T_299 <= 58'h0;
    end else if (csr_wen) begin
      if (_T_998) begin
        _T_299 <= wdata[63:6];
      end else if (_T_297[6]) begin
        _T_299 <= _T_302;
      end
    end else if (_T_297[6]) begin
      _T_299 <= _T_302;
    end
  end
  always @(posedge clock) begin
    if(CSRFile_cov_write_en & CSRFile_cov_write_mask) begin
      CSRFile_cov[CSRFile_cov_write_addr] <= CSRFile_cov_write_data; // @[Coverage map for CSRFile]
    end
  end
endmodule
module BreakpointUnit(
  input         io_status_debug,
  input  [1:0]  io_status_prv,
  input         io_bp_0_control_action,
  input  [1:0]  io_bp_0_control_tmatch,
  input         io_bp_0_control_m,
  input         io_bp_0_control_s,
  input         io_bp_0_control_u,
  input         io_bp_0_control_x,
  input         io_bp_0_control_w,
  input         io_bp_0_control_r,
  input  [38:0] io_bp_0_address,
  input  [38:0] io_pc,
  input  [38:0] io_ea,
  output        io_xcpt_if,
  output        io_xcpt_ld,
  output        io_xcpt_st,
  output        io_debug_if,
  output        io_debug_ld,
  output        io_debug_st,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [3:0] _T_22; // @[Cat.scala 30:58]
  wire [3:0] _T_23; // @[Breakpoint.scala 30:68]
  wire  _T_25; // @[Breakpoint.scala 30:50]
  wire  _T_27; // @[Breakpoint.scala 73:22]
  wire  _T_29; // @[Breakpoint.scala 44:8]
  wire  _T_31; // @[Breakpoint.scala 44:20]
  wire  _T_35; // @[Breakpoint.scala 38:73]
  wire  _T_37; // @[Breakpoint.scala 38:73]
  wire  _T_39; // @[Breakpoint.scala 38:73]
  wire [3:0] _T_42; // @[Cat.scala 30:58]
  wire [38:0] _GEN_6; // @[Breakpoint.scala 41:9]
  wire [38:0] _T_43; // @[Breakpoint.scala 41:9]
  wire [38:0] _T_55; // @[Breakpoint.scala 41:33]
  wire  _T_56; // @[Breakpoint.scala 41:19]
  wire  _T_57; // @[Breakpoint.scala 47:8]
  wire  _T_58; // @[Breakpoint.scala 73:38]
  wire  _T_60; // @[Breakpoint.scala 74:22]
  wire  _T_91; // @[Breakpoint.scala 74:38]
  wire  _T_93; // @[Breakpoint.scala 75:22]
  wire  _T_95; // @[Breakpoint.scala 44:8]
  wire  _T_97; // @[Breakpoint.scala 44:20]
  wire [38:0] _T_109; // @[Breakpoint.scala 41:9]
  wire  _T_122; // @[Breakpoint.scala 41:19]
  wire  _T_123; // @[Breakpoint.scala 47:8]
  wire  _T_124; // @[Breakpoint.scala 75:38]
  wire [29:0] BreakpointUnit_covSum;
  assign _T_22 = {io_bp_0_control_m,1'h0,io_bp_0_control_s,io_bp_0_control_u}; // @[Cat.scala 30:58]
  assign _T_23 = _T_22 >> io_status_prv; // @[Breakpoint.scala 30:68]
  assign _T_25 = ~io_status_debug & _T_23[0]; // @[Breakpoint.scala 30:50]
  assign _T_27 = _T_25 & io_bp_0_control_r; // @[Breakpoint.scala 73:22]
  assign _T_29 = io_ea >= io_bp_0_address; // @[Breakpoint.scala 44:8]
  assign _T_31 = _T_29 ^ io_bp_0_control_tmatch[0]; // @[Breakpoint.scala 44:20]
  assign _T_35 = io_bp_0_control_tmatch[0] & io_bp_0_address[0]; // @[Breakpoint.scala 38:73]
  assign _T_37 = _T_35 & io_bp_0_address[1]; // @[Breakpoint.scala 38:73]
  assign _T_39 = _T_37 & io_bp_0_address[2]; // @[Breakpoint.scala 38:73]
  assign _T_42 = {_T_39,_T_37,_T_35,io_bp_0_control_tmatch[0]}; // @[Cat.scala 30:58]
  assign _GEN_6 = {{35'd0}, _T_42}; // @[Breakpoint.scala 41:9]
  assign _T_43 = ~io_ea | _GEN_6; // @[Breakpoint.scala 41:9]
  assign _T_55 = ~io_bp_0_address | _GEN_6; // @[Breakpoint.scala 41:33]
  assign _T_56 = _T_43 == _T_55; // @[Breakpoint.scala 41:19]
  assign _T_57 = io_bp_0_control_tmatch[1] ? _T_31 : _T_56; // @[Breakpoint.scala 47:8]
  assign _T_58 = _T_27 & _T_57; // @[Breakpoint.scala 73:38]
  assign _T_60 = _T_25 & io_bp_0_control_w; // @[Breakpoint.scala 74:22]
  assign _T_91 = _T_60 & _T_57; // @[Breakpoint.scala 74:38]
  assign _T_93 = _T_25 & io_bp_0_control_x; // @[Breakpoint.scala 75:22]
  assign _T_95 = io_pc >= io_bp_0_address; // @[Breakpoint.scala 44:8]
  assign _T_97 = _T_95 ^ io_bp_0_control_tmatch[0]; // @[Breakpoint.scala 44:20]
  assign _T_109 = ~io_pc | _GEN_6; // @[Breakpoint.scala 41:9]
  assign _T_122 = _T_109 == _T_55; // @[Breakpoint.scala 41:19]
  assign _T_123 = io_bp_0_control_tmatch[1] ? _T_97 : _T_122; // @[Breakpoint.scala 47:8]
  assign _T_124 = _T_93 & _T_123; // @[Breakpoint.scala 75:38]
  assign io_xcpt_if = _T_124 & ~io_bp_0_control_action; // @[Breakpoint.scala 64:14 Breakpoint.scala 80:34]
  assign io_xcpt_ld = _T_58 & ~io_bp_0_control_action; // @[Breakpoint.scala 65:14 Breakpoint.scala 78:34]
  assign io_xcpt_st = _T_91 & ~io_bp_0_control_action; // @[Breakpoint.scala 66:14 Breakpoint.scala 79:34]
  assign io_debug_if = _T_124 & io_bp_0_control_action; // @[Breakpoint.scala 67:15 Breakpoint.scala 80:69]
  assign io_debug_ld = _T_58 & io_bp_0_control_action; // @[Breakpoint.scala 68:15 Breakpoint.scala 78:69]
  assign io_debug_st = _T_91 & io_bp_0_control_action; // @[Breakpoint.scala 69:15 Breakpoint.scala 79:69]
  assign BreakpointUnit_covSum = 30'h0;
  assign io_covSum = BreakpointUnit_covSum;
  assign metaAssert = 1'h0;
endmodule
module ALU(
  input         io_dw,
  input  [3:0]  io_fn,
  input  [63:0] io_in2,
  input  [63:0] io_in1,
  output [63:0] io_out,
  output [63:0] io_adder_out,
  output        io_cmp_out,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [63:0] in2_inv; // @[ALU.scala 62:20]
  wire [63:0] in1_xor_in2; // @[ALU.scala 63:28]
  wire [63:0] _T_14; // @[ALU.scala 64:26]
  wire [63:0] _GEN_1; // @[ALU.scala 64:36]
  wire  _T_20; // @[ALU.scala 68:24]
  wire  _T_25; // @[ALU.scala 69:8]
  wire  slt; // @[ALU.scala 68:8]
  wire  _T_29; // @[ALU.scala 70:68]
  wire  _T_30; // @[ALU.scala 70:41]
  wire  _T_34; // @[ALU.scala 77:46]
  wire [31:0] _T_36; // @[Bitwise.scala 72:12]
  wire [31:0] _T_39; // @[ALU.scala 78:24]
  wire  _T_42; // @[ALU.scala 79:33]
  wire [5:0] shamt; // @[Cat.scala 30:58]
  wire [63:0] shin_r; // @[Cat.scala 30:58]
  wire  _T_45; // @[ALU.scala 82:24]
  wire  _T_46; // @[ALU.scala 82:44]
  wire  _T_47; // @[ALU.scala 82:35]
  wire [63:0] _T_51; // @[Bitwise.scala 103:31]
  wire [63:0] _T_53; // @[Bitwise.scala 103:65]
  wire [63:0] _T_55; // @[Bitwise.scala 103:75]
  wire [63:0] _T_56; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_2; // @[Bitwise.scala 103:31]
  wire [63:0] _T_61; // @[Bitwise.scala 103:31]
  wire [63:0] _T_63; // @[Bitwise.scala 103:65]
  wire [63:0] _T_65; // @[Bitwise.scala 103:75]
  wire [63:0] _T_66; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_3; // @[Bitwise.scala 103:31]
  wire [63:0] _T_71; // @[Bitwise.scala 103:31]
  wire [63:0] _T_73; // @[Bitwise.scala 103:65]
  wire [63:0] _T_75; // @[Bitwise.scala 103:75]
  wire [63:0] _T_76; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_4; // @[Bitwise.scala 103:31]
  wire [63:0] _T_81; // @[Bitwise.scala 103:31]
  wire [63:0] _T_83; // @[Bitwise.scala 103:65]
  wire [63:0] _T_85; // @[Bitwise.scala 103:75]
  wire [63:0] _T_86; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_5; // @[Bitwise.scala 103:31]
  wire [63:0] _T_91; // @[Bitwise.scala 103:31]
  wire [63:0] _T_93; // @[Bitwise.scala 103:65]
  wire [63:0] _T_95; // @[Bitwise.scala 103:75]
  wire [63:0] _T_96; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_6; // @[Bitwise.scala 103:31]
  wire [63:0] _T_101; // @[Bitwise.scala 103:31]
  wire [63:0] _T_103; // @[Bitwise.scala 103:65]
  wire [63:0] _T_105; // @[Bitwise.scala 103:75]
  wire [63:0] _T_106; // @[Bitwise.scala 103:39]
  wire [63:0] shin; // @[ALU.scala 82:17]
  wire  _T_109; // @[ALU.scala 83:35]
  wire [64:0] _T_111; // @[ALU.scala 83:57]
  wire [64:0] _T_112; // @[ALU.scala 83:64]
  wire [63:0] shout_r; // @[ALU.scala 83:73]
  wire [63:0] _T_116; // @[Bitwise.scala 103:31]
  wire [63:0] _T_118; // @[Bitwise.scala 103:65]
  wire [63:0] _T_120; // @[Bitwise.scala 103:75]
  wire [63:0] _T_121; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_7; // @[Bitwise.scala 103:31]
  wire [63:0] _T_126; // @[Bitwise.scala 103:31]
  wire [63:0] _T_128; // @[Bitwise.scala 103:65]
  wire [63:0] _T_130; // @[Bitwise.scala 103:75]
  wire [63:0] _T_131; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_8; // @[Bitwise.scala 103:31]
  wire [63:0] _T_136; // @[Bitwise.scala 103:31]
  wire [63:0] _T_138; // @[Bitwise.scala 103:65]
  wire [63:0] _T_140; // @[Bitwise.scala 103:75]
  wire [63:0] _T_141; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_9; // @[Bitwise.scala 103:31]
  wire [63:0] _T_146; // @[Bitwise.scala 103:31]
  wire [63:0] _T_148; // @[Bitwise.scala 103:65]
  wire [63:0] _T_150; // @[Bitwise.scala 103:75]
  wire [63:0] _T_151; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_10; // @[Bitwise.scala 103:31]
  wire [63:0] _T_156; // @[Bitwise.scala 103:31]
  wire [63:0] _T_158; // @[Bitwise.scala 103:65]
  wire [63:0] _T_160; // @[Bitwise.scala 103:75]
  wire [63:0] _T_161; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_11; // @[Bitwise.scala 103:31]
  wire [63:0] _T_166; // @[Bitwise.scala 103:31]
  wire [63:0] _T_168; // @[Bitwise.scala 103:65]
  wire [63:0] _T_170; // @[Bitwise.scala 103:75]
  wire [63:0] shout_l; // @[Bitwise.scala 103:39]
  wire [63:0] _T_174; // @[ALU.scala 85:18]
  wire  _T_175; // @[ALU.scala 86:25]
  wire [63:0] _T_176; // @[ALU.scala 86:18]
  wire [63:0] shout; // @[ALU.scala 85:74]
  wire  _T_177; // @[ALU.scala 89:25]
  wire  _T_178; // @[ALU.scala 89:45]
  wire  _T_179; // @[ALU.scala 89:36]
  wire [63:0] _T_180; // @[ALU.scala 89:18]
  wire  _T_182; // @[ALU.scala 90:44]
  wire  _T_183; // @[ALU.scala 90:35]
  wire [63:0] _T_184; // @[ALU.scala 90:63]
  wire [63:0] _T_185; // @[ALU.scala 90:18]
  wire [63:0] logic_; // @[ALU.scala 89:78]
  wire  _T_186; // @[ALU.scala 41:30]
  wire  _T_187; // @[ALU.scala 91:35]
  wire [63:0] _GEN_12; // @[ALU.scala 91:43]
  wire [63:0] _T_188; // @[ALU.scala 91:43]
  wire [63:0] shift_logic; // @[ALU.scala 91:51]
  wire  _T_189; // @[ALU.scala 92:23]
  wire  _T_190; // @[ALU.scala 92:43]
  wire  _T_191; // @[ALU.scala 92:34]
  wire [63:0] out; // @[ALU.scala 92:16]
  wire [31:0] _T_195; // @[Bitwise.scala 72:12]
  wire [63:0] _T_197; // @[Cat.scala 30:58]
  wire [29:0] ALU_covSum;
  assign in2_inv = io_fn[3] ? ~io_in2 : io_in2; // @[ALU.scala 62:20]
  assign in1_xor_in2 = io_in1 ^ in2_inv; // @[ALU.scala 63:28]
  assign _T_14 = io_in1 + in2_inv; // @[ALU.scala 64:26]
  assign _GEN_1 = {{63'd0}, io_fn[3]}; // @[ALU.scala 64:36]
  assign _T_20 = io_in1[63] == io_in2[63]; // @[ALU.scala 68:24]
  assign _T_25 = io_fn[1] ? io_in2[63] : io_in1[63]; // @[ALU.scala 69:8]
  assign slt = _T_20 ? io_adder_out[63] : _T_25; // @[ALU.scala 68:8]
  assign _T_29 = in1_xor_in2 == 64'h0; // @[ALU.scala 70:68]
  assign _T_30 = io_fn[3] ? slt : _T_29; // @[ALU.scala 70:41]
  assign _T_34 = io_fn[3] & io_in1[31]; // @[ALU.scala 77:46]
  assign _T_36 = _T_34 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  assign _T_39 = io_dw ? io_in1[63:32] : _T_36; // @[ALU.scala 78:24]
  assign _T_42 = io_in2[5] & io_dw; // @[ALU.scala 79:33]
  assign shamt = {_T_42,io_in2[4:0]}; // @[Cat.scala 30:58]
  assign shin_r = {_T_39,io_in1[31:0]}; // @[Cat.scala 30:58]
  assign _T_45 = io_fn == 4'h5; // @[ALU.scala 82:24]
  assign _T_46 = io_fn == 4'hb; // @[ALU.scala 82:44]
  assign _T_47 = _T_45 | _T_46; // @[ALU.scala 82:35]
  assign _T_51 = {{32'd0}, shin_r[63:32]}; // @[Bitwise.scala 103:31]
  assign _T_53 = {shin_r[31:0], 32'h0}; // @[Bitwise.scala 103:65]
  assign _T_55 = _T_53 & 64'hffffffff00000000; // @[Bitwise.scala 103:75]
  assign _T_56 = _T_51 | _T_55; // @[Bitwise.scala 103:39]
  assign _GEN_2 = {{16'd0}, _T_56[63:16]}; // @[Bitwise.scala 103:31]
  assign _T_61 = _GEN_2 & 64'hffff0000ffff; // @[Bitwise.scala 103:31]
  assign _T_63 = {_T_56[47:0], 16'h0}; // @[Bitwise.scala 103:65]
  assign _T_65 = _T_63 & 64'hffff0000ffff0000; // @[Bitwise.scala 103:75]
  assign _T_66 = _T_61 | _T_65; // @[Bitwise.scala 103:39]
  assign _GEN_3 = {{8'd0}, _T_66[63:8]}; // @[Bitwise.scala 103:31]
  assign _T_71 = _GEN_3 & 64'hff00ff00ff00ff; // @[Bitwise.scala 103:31]
  assign _T_73 = {_T_66[55:0], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_75 = _T_73 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 103:75]
  assign _T_76 = _T_71 | _T_75; // @[Bitwise.scala 103:39]
  assign _GEN_4 = {{4'd0}, _T_76[63:4]}; // @[Bitwise.scala 103:31]
  assign _T_81 = _GEN_4 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 103:31]
  assign _T_83 = {_T_76[59:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_85 = _T_83 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 103:75]
  assign _T_86 = _T_81 | _T_85; // @[Bitwise.scala 103:39]
  assign _GEN_5 = {{2'd0}, _T_86[63:2]}; // @[Bitwise.scala 103:31]
  assign _T_91 = _GEN_5 & 64'h3333333333333333; // @[Bitwise.scala 103:31]
  assign _T_93 = {_T_86[61:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_95 = _T_93 & 64'hcccccccccccccccc; // @[Bitwise.scala 103:75]
  assign _T_96 = _T_91 | _T_95; // @[Bitwise.scala 103:39]
  assign _GEN_6 = {{1'd0}, _T_96[63:1]}; // @[Bitwise.scala 103:31]
  assign _T_101 = _GEN_6 & 64'h5555555555555555; // @[Bitwise.scala 103:31]
  assign _T_103 = {_T_96[62:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_105 = _T_103 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 103:75]
  assign _T_106 = _T_101 | _T_105; // @[Bitwise.scala 103:39]
  assign shin = _T_47 ? shin_r : _T_106; // @[ALU.scala 82:17]
  assign _T_109 = io_fn[3] & shin[63]; // @[ALU.scala 83:35]
  assign _T_111 = {_T_109,shin}; // @[ALU.scala 83:57]
  assign _T_112 = $signed(_T_111) >>> shamt; // @[ALU.scala 83:64]
  assign shout_r = _T_112[63:0]; // @[ALU.scala 83:73]
  assign _T_116 = {{32'd0}, shout_r[63:32]}; // @[Bitwise.scala 103:31]
  assign _T_118 = {shout_r[31:0], 32'h0}; // @[Bitwise.scala 103:65]
  assign _T_120 = _T_118 & 64'hffffffff00000000; // @[Bitwise.scala 103:75]
  assign _T_121 = _T_116 | _T_120; // @[Bitwise.scala 103:39]
  assign _GEN_7 = {{16'd0}, _T_121[63:16]}; // @[Bitwise.scala 103:31]
  assign _T_126 = _GEN_7 & 64'hffff0000ffff; // @[Bitwise.scala 103:31]
  assign _T_128 = {_T_121[47:0], 16'h0}; // @[Bitwise.scala 103:65]
  assign _T_130 = _T_128 & 64'hffff0000ffff0000; // @[Bitwise.scala 103:75]
  assign _T_131 = _T_126 | _T_130; // @[Bitwise.scala 103:39]
  assign _GEN_8 = {{8'd0}, _T_131[63:8]}; // @[Bitwise.scala 103:31]
  assign _T_136 = _GEN_8 & 64'hff00ff00ff00ff; // @[Bitwise.scala 103:31]
  assign _T_138 = {_T_131[55:0], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_140 = _T_138 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 103:75]
  assign _T_141 = _T_136 | _T_140; // @[Bitwise.scala 103:39]
  assign _GEN_9 = {{4'd0}, _T_141[63:4]}; // @[Bitwise.scala 103:31]
  assign _T_146 = _GEN_9 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 103:31]
  assign _T_148 = {_T_141[59:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_150 = _T_148 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 103:75]
  assign _T_151 = _T_146 | _T_150; // @[Bitwise.scala 103:39]
  assign _GEN_10 = {{2'd0}, _T_151[63:2]}; // @[Bitwise.scala 103:31]
  assign _T_156 = _GEN_10 & 64'h3333333333333333; // @[Bitwise.scala 103:31]
  assign _T_158 = {_T_151[61:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_160 = _T_158 & 64'hcccccccccccccccc; // @[Bitwise.scala 103:75]
  assign _T_161 = _T_156 | _T_160; // @[Bitwise.scala 103:39]
  assign _GEN_11 = {{1'd0}, _T_161[63:1]}; // @[Bitwise.scala 103:31]
  assign _T_166 = _GEN_11 & 64'h5555555555555555; // @[Bitwise.scala 103:31]
  assign _T_168 = {_T_161[62:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_170 = _T_168 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 103:75]
  assign shout_l = _T_166 | _T_170; // @[Bitwise.scala 103:39]
  assign _T_174 = _T_47 ? shout_r : 64'h0; // @[ALU.scala 85:18]
  assign _T_175 = io_fn == 4'h1; // @[ALU.scala 86:25]
  assign _T_176 = _T_175 ? shout_l : 64'h0; // @[ALU.scala 86:18]
  assign shout = _T_174 | _T_176; // @[ALU.scala 85:74]
  assign _T_177 = io_fn == 4'h4; // @[ALU.scala 89:25]
  assign _T_178 = io_fn == 4'h6; // @[ALU.scala 89:45]
  assign _T_179 = _T_177 | _T_178; // @[ALU.scala 89:36]
  assign _T_180 = _T_179 ? in1_xor_in2 : 64'h0; // @[ALU.scala 89:18]
  assign _T_182 = io_fn == 4'h7; // @[ALU.scala 90:44]
  assign _T_183 = _T_178 | _T_182; // @[ALU.scala 90:35]
  assign _T_184 = io_in1 & io_in2; // @[ALU.scala 90:63]
  assign _T_185 = _T_183 ? _T_184 : 64'h0; // @[ALU.scala 90:18]
  assign logic_ = _T_180 | _T_185; // @[ALU.scala 89:78]
  assign _T_186 = io_fn >= 4'hc; // @[ALU.scala 41:30]
  assign _T_187 = _T_186 & slt; // @[ALU.scala 91:35]
  assign _GEN_12 = {{63'd0}, _T_187}; // @[ALU.scala 91:43]
  assign _T_188 = _GEN_12 | logic_; // @[ALU.scala 91:43]
  assign shift_logic = _T_188 | shout; // @[ALU.scala 91:51]
  assign _T_189 = io_fn == 4'h0; // @[ALU.scala 92:23]
  assign _T_190 = io_fn == 4'ha; // @[ALU.scala 92:43]
  assign _T_191 = _T_189 | _T_190; // @[ALU.scala 92:34]
  assign out = _T_191 ? io_adder_out : shift_logic; // @[ALU.scala 92:16]
  assign _T_195 = out[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  assign _T_197 = {_T_195,out[31:0]}; // @[Cat.scala 30:58]
  assign io_out = io_dw ? out : _T_197; // @[ALU.scala 94:10 ALU.scala 97:37]
  assign io_adder_out = _T_14 + _GEN_1; // @[ALU.scala 64:16]
  assign io_cmp_out = io_fn[0] ^ _T_30; // @[ALU.scala 70:14]
  assign ALU_covSum = 30'h0;
  assign io_covSum = ALU_covSum;
  assign metaAssert = 1'h0;
endmodule
module MulDiv(
  input         clock,
  input         reset,
  output        io_req_ready,
  input         io_req_valid,
  input  [3:0]  io_req_bits_fn,
  input         io_req_bits_dw,
  input  [63:0] io_req_bits_in1,
  input  [63:0] io_req_bits_in2,
  input  [4:0]  io_req_bits_tag,
  input         io_kill,
  input         io_resp_ready,
  output        io_resp_valid,
  output [63:0] io_resp_bits_data,
  output [4:0]  io_resp_bits_tag,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [2:0] state; // @[Multiplier.scala 51:18]
  reg [31:0] _RAND_0;
  reg  req_dw; // @[Multiplier.scala 53:16]
  reg [31:0] _RAND_1;
  reg [4:0] req_tag; // @[Multiplier.scala 53:16]
  reg [31:0] _RAND_2;
  reg [6:0] count; // @[Multiplier.scala 54:18]
  reg [31:0] _RAND_3;
  reg  neg_out; // @[Multiplier.scala 57:20]
  reg [31:0] _RAND_4;
  reg  isHi; // @[Multiplier.scala 58:17]
  reg [31:0] _RAND_5;
  reg  resHi; // @[Multiplier.scala 59:18]
  reg [31:0] _RAND_6;
  reg [64:0] divisor; // @[Multiplier.scala 60:20]
  reg [95:0] _RAND_7;
  reg [129:0] remainder; // @[Multiplier.scala 61:22]
  reg [159:0] _RAND_8;
  wire [3:0] _T_22; // @[Decode.scala 14:65]
  wire  cmdMul; // @[Decode.scala 14:121]
  wire [3:0] _T_25; // @[Decode.scala 14:65]
  wire  _T_26; // @[Decode.scala 14:121]
  wire [3:0] _T_27; // @[Decode.scala 14:65]
  wire  _T_28; // @[Decode.scala 14:121]
  wire  cmdHi; // @[Decode.scala 15:30]
  wire [3:0] _T_31; // @[Decode.scala 14:65]
  wire  _T_32; // @[Decode.scala 14:121]
  wire [3:0] _T_33; // @[Decode.scala 14:65]
  wire  _T_34; // @[Decode.scala 14:121]
  wire  lhsSigned; // @[Decode.scala 15:30]
  wire  _T_38; // @[Decode.scala 14:121]
  wire  rhsSigned; // @[Decode.scala 15:30]
  wire  _T_45; // @[Multiplier.scala 81:29]
  wire  lhs_sign; // @[Multiplier.scala 81:23]
  wire [31:0] _T_47; // @[Bitwise.scala 72:12]
  wire [31:0] _T_49; // @[Multiplier.scala 82:17]
  wire [63:0] lhs_in; // @[Cat.scala 30:58]
  wire  _T_55; // @[Multiplier.scala 81:29]
  wire  rhs_sign; // @[Multiplier.scala 81:23]
  wire [31:0] _T_57; // @[Bitwise.scala 72:12]
  wire [31:0] _T_59; // @[Multiplier.scala 82:17]
  wire [64:0] subtractor; // @[Multiplier.scala 88:37]
  wire [63:0] result; // @[Multiplier.scala 89:19]
  wire [63:0] negated_remainder; // @[Multiplier.scala 90:27]
  wire  _T_68; // @[Multiplier.scala 92:39]
  wire  _T_71; // @[Multiplier.scala 101:39]
  wire  _T_72; // @[Multiplier.scala 106:39]
  wire [128:0] _T_75; // @[Cat.scala 30:58]
  wire [64:0] _T_79; // @[Multiplier.scala 110:37]
  wire [8:0] _T_83; // @[Multiplier.scala 112:60]
  wire [64:0] _GEN_37; // @[Multiplier.scala 112:67]
  wire [73:0] _T_84; // @[Multiplier.scala 112:67]
  wire [73:0] _GEN_38; // @[Multiplier.scala 112:76]
  wire [73:0] _T_89; // @[Cat.scala 30:58]
  wire [129:0] _T_90; // @[Cat.scala 30:58]
  wire  _T_91; // @[Multiplier.scala 114:32]
  wire  _T_92; // @[Multiplier.scala 114:57]
  wire [10:0] _T_93; // @[Multiplier.scala 116:56]
  wire [64:0] _T_95; // @[Multiplier.scala 116:46]
  wire  _T_97; // @[Multiplier.scala 117:47]
  wire  _T_99; // @[Multiplier.scala 117:81]
  wire  _T_100; // @[Multiplier.scala 117:72]
  wire  _T_102; // @[Multiplier.scala 117:87]
  wire [63:0] _T_104; // @[Multiplier.scala 118:24]
  wire  _T_105; // @[Multiplier.scala 118:37]
  wire  _T_106; // @[Multiplier.scala 118:13]
  wire [10:0] _T_110; // @[Multiplier.scala 119:36]
  wire [128:0] _T_112; // @[Multiplier.scala 119:27]
  wire [129:0] _T_114; // @[Multiplier.scala 120:55]
  wire [128:0] _T_116; // @[Cat.scala 30:58]
  wire [129:0] _T_120; // @[Cat.scala 30:58]
  wire [6:0] _T_122; // @[Multiplier.scala 123:20]
  wire  _T_123; // @[Multiplier.scala 124:25]
  wire  _T_124; // @[Multiplier.scala 124:16]
  wire  _T_125; // @[Multiplier.scala 129:39]
  wire [63:0] _T_129; // @[Multiplier.scala 134:14]
  wire [128:0] _T_133; // @[Cat.scala 30:58]
  wire  _T_134; // @[Multiplier.scala 138:17]
  wire  _T_138; // @[Multiplier.scala 146:24]
  wire  _T_141; // @[Multiplier.scala 146:30]
  wire  _T_146; // @[CircuitMath.scala 37:22]
  wire  _T_149; // @[CircuitMath.scala 37:22]
  wire  _T_152; // @[CircuitMath.scala 37:22]
  wire  _T_155; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_159; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_160; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_164; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_165; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_166; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_167; // @[Cat.scala 30:58]
  wire  _T_170; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_174; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_175; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_179; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_180; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_181; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_182; // @[Cat.scala 30:58]
  wire [2:0] _T_183; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_184; // @[Cat.scala 30:58]
  wire  _T_187; // @[CircuitMath.scala 37:22]
  wire  _T_190; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_194; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_195; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_199; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_200; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_201; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_202; // @[Cat.scala 30:58]
  wire  _T_205; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_209; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_210; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_214; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_215; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_216; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_217; // @[Cat.scala 30:58]
  wire [2:0] _T_218; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_219; // @[Cat.scala 30:58]
  wire [3:0] _T_220; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_221; // @[Cat.scala 30:58]
  wire  _T_224; // @[CircuitMath.scala 37:22]
  wire  _T_227; // @[CircuitMath.scala 37:22]
  wire  _T_230; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_234; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_235; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_239; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_240; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_241; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_242; // @[Cat.scala 30:58]
  wire  _T_245; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_249; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_250; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_254; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_255; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_256; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_257; // @[Cat.scala 30:58]
  wire [2:0] _T_258; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_259; // @[Cat.scala 30:58]
  wire  _T_262; // @[CircuitMath.scala 37:22]
  wire  _T_265; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_269; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_270; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_274; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_275; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_276; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_277; // @[Cat.scala 30:58]
  wire  _T_280; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_284; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_285; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_289; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_290; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_291; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_292; // @[Cat.scala 30:58]
  wire [2:0] _T_293; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_294; // @[Cat.scala 30:58]
  wire [3:0] _T_295; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_296; // @[Cat.scala 30:58]
  wire [4:0] _T_297; // @[CircuitMath.scala 38:21]
  wire [5:0] _T_298; // @[Cat.scala 30:58]
  wire  _T_303; // @[CircuitMath.scala 37:22]
  wire  _T_306; // @[CircuitMath.scala 37:22]
  wire  _T_309; // @[CircuitMath.scala 37:22]
  wire  _T_312; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_316; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_317; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_321; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_322; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_323; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_324; // @[Cat.scala 30:58]
  wire  _T_327; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_331; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_332; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_336; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_337; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_338; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_339; // @[Cat.scala 30:58]
  wire [2:0] _T_340; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_341; // @[Cat.scala 30:58]
  wire  _T_344; // @[CircuitMath.scala 37:22]
  wire  _T_347; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_351; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_352; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_356; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_357; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_358; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_359; // @[Cat.scala 30:58]
  wire  _T_362; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_366; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_367; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_371; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_372; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_373; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_374; // @[Cat.scala 30:58]
  wire [2:0] _T_375; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_376; // @[Cat.scala 30:58]
  wire [3:0] _T_377; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_378; // @[Cat.scala 30:58]
  wire  _T_381; // @[CircuitMath.scala 37:22]
  wire  _T_384; // @[CircuitMath.scala 37:22]
  wire  _T_387; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_391; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_392; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_396; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_397; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_398; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_399; // @[Cat.scala 30:58]
  wire  _T_402; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_406; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_407; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_411; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_412; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_413; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_414; // @[Cat.scala 30:58]
  wire [2:0] _T_415; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_416; // @[Cat.scala 30:58]
  wire  _T_419; // @[CircuitMath.scala 37:22]
  wire  _T_422; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_426; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_427; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_431; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_432; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_433; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_434; // @[Cat.scala 30:58]
  wire  _T_437; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_441; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_442; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_446; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_447; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_448; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_449; // @[Cat.scala 30:58]
  wire [2:0] _T_450; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_451; // @[Cat.scala 30:58]
  wire [3:0] _T_452; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_453; // @[Cat.scala 30:58]
  wire [4:0] _T_454; // @[CircuitMath.scala 38:21]
  wire [5:0] _T_455; // @[Cat.scala 30:58]
  wire [5:0] _T_460; // @[Multiplier.scala 152:35]
  wire  _T_464; // @[Multiplier.scala 153:30]
  wire  _T_465; // @[Multiplier.scala 153:52]
  wire  _T_466; // @[Multiplier.scala 153:41]
  wire [126:0] _GEN_39; // @[Multiplier.scala 155:39]
  wire [126:0] _T_468; // @[Multiplier.scala 155:39]
  wire [128:0] _GEN_16; // @[Multiplier.scala 154:19]
  wire  _T_471; // @[Multiplier.scala 159:18]
  wire  _T_472; // @[Decoupled.scala 37:37]
  wire  _T_473; // @[Multiplier.scala 161:24]
  wire  _T_474; // @[Decoupled.scala 37:37]
  wire  _T_475; // @[Multiplier.scala 165:46]
  wire  _T_480; // @[Multiplier.scala 168:46]
  wire [2:0] _T_481; // @[Multiplier.scala 168:38]
  wire  _T_482; // @[Multiplier.scala 169:46]
  wire [64:0] _T_484; // @[Cat.scala 30:58]
  wire [2:0] _T_486; // @[Multiplier.scala 175:23]
  wire  outMul; // @[Multiplier.scala 175:52]
  wire  _T_492; // @[Multiplier.scala 176:52]
  wire [31:0] loOut; // @[Multiplier.scala 176:18]
  wire [31:0] _T_499; // @[Bitwise.scala 72:12]
  wire [31:0] hiOut; // @[Multiplier.scala 177:18]
  wire  _T_502; // @[Multiplier.scala 180:27]
  wire  _T_503; // @[Multiplier.scala 180:51]
  reg [19:0] MulDiv_state; // @[Register tracking MulDiv state]
  reg [31:0] _RAND_9;
  reg  MulDiv_cov [0:1048575]; // @[Coverage map for MulDiv]
  reg [31:0] _RAND_10;
  wire  MulDiv_cov_read_data; // @[Coverage map for MulDiv]
  wire [19:0] MulDiv_cov_read_addr; // @[Coverage map for MulDiv]
  wire  MulDiv_cov_write_data; // @[Coverage map for MulDiv]
  wire [19:0] MulDiv_cov_write_addr; // @[Coverage map for MulDiv]
  wire  MulDiv_cov_write_mask; // @[Coverage map for MulDiv]
  wire  MulDiv_cov_write_en; // @[Coverage map for MulDiv]
  reg [29:0] MulDiv_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_11;
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  mux_cond_4;
  wire  mux_cond_5;
  wire  mux_cond_6;
  wire  mux_cond_7;
  wire  mux_cond_8;
  wire  mux_cond_9;
  wire  mux_cond_10;
  wire  mux_cond_11;
  wire  mux_cond_12;
  wire  mux_cond_13;
  wire  mux_cond_14;
  wire  mux_cond_15;
  wire  mux_cond_16;
  wire  mux_cond_17;
  wire  mux_cond_18;
  wire  mux_cond_19;
  wire  mux_cond_20;
  wire  mux_cond_21;
  wire  mux_cond_22;
  wire  mux_cond_23;
  wire  mux_cond_24;
  wire  mux_cond_25;
  wire  mux_cond_26;
  wire  mux_cond_27;
  wire  mux_cond_28;
  wire  mux_cond_29;
  wire  mux_cond_30;
  wire  mux_cond_31;
  wire  mux_cond_32;
  wire  mux_cond_33;
  wire  mux_cond_34;
  wire  mux_cond_35;
  wire  mux_cond_36;
  wire  mux_cond_37;
  wire  mux_cond_38;
  wire  mux_cond_39;
  wire  mux_cond_40;
  wire  mux_cond_41;
  wire  mux_cond_42;
  wire  mux_cond_43;
  wire  mux_cond_44;
  wire  mux_cond_45;
  wire  mux_cond_46;
  wire  mux_cond_47;
  wire  mux_cond_48;
  wire  mux_cond_49;
  wire  mux_cond_50;
  wire  mux_cond_51;
  wire  mux_cond_52;
  wire  mux_cond_53;
  wire  mux_cond_54;
  wire  mux_cond_55;
  wire  mux_cond_56;
  wire  mux_cond_57;
  wire  mux_cond_58;
  wire  mux_cond_59;
  wire  mux_cond_60;
  wire  mux_cond_61;
  wire  mux_cond_62;
  wire  mux_cond_63;
  wire  mux_cond_64;
  wire  mux_cond_65;
  wire  mux_cond_66;
  wire  mux_cond_67;
  wire  mux_cond_68;
  wire  mux_cond_69;
  wire  mux_cond_70;
  wire  mux_cond_71;
  wire  mux_cond_72;
  wire  mux_cond_73;
  wire  mux_cond_74;
  wire  mux_cond_75;
  wire  mux_cond_76;
  wire  mux_cond_77;
  wire  mux_cond_78;
  wire  mux_cond_79;
  wire  mux_cond_80;
  wire  mux_cond_81;
  wire  mux_cond_82;
  wire  mux_cond_83;
  wire  mux_cond_84;
  wire  mux_cond_85;
  wire  mux_cond_86;
  wire  mux_cond_87;
  wire  mux_cond_88;
  wire  mux_cond_89;
  wire  mux_cond_90;
  wire  mux_cond_91;
  wire  mux_cond_92;
  wire  mux_cond_93;
  wire  mux_cond_94;
  wire  mux_cond_95;
  wire  mux_cond_96;
  wire  mux_cond_97;
  wire [10:0] resHi_shl;
  wire [19:0] resHi_pad;
  wire [13:0] state_shl;
  wire [19:0] state_pad;
  wire [5:0] req_dw_shl;
  wire [19:0] req_dw_pad;
  wire [16:0] neg_out_shl;
  wire [19:0] neg_out_pad;
  wire [13:0] isHi_shl;
  wire [19:0] isHi_pad;
  wire [8:0] mux_cond_0_shl;
  wire [19:0] mux_cond_0_pad;
  wire  mux_cond_1_shl;
  wire [19:0] mux_cond_1_pad;
  wire [11:0] mux_cond_2_shl;
  wire [19:0] mux_cond_2_pad;
  wire [9:0] mux_cond_3_shl;
  wire [19:0] mux_cond_3_pad;
  wire [7:0] mux_cond_4_shl;
  wire [19:0] mux_cond_4_pad;
  wire [5:0] mux_cond_5_shl;
  wire [19:0] mux_cond_5_pad;
  wire [12:0] mux_cond_6_shl;
  wire [19:0] mux_cond_6_pad;
  wire [9:0] mux_cond_7_shl;
  wire [19:0] mux_cond_7_pad;
  wire [2:0] mux_cond_8_shl;
  wire [19:0] mux_cond_8_pad;
  wire [1:0] mux_cond_9_shl;
  wire [19:0] mux_cond_9_pad;
  wire [12:0] mux_cond_10_shl;
  wire [19:0] mux_cond_10_pad;
  wire [8:0] mux_cond_11_shl;
  wire [19:0] mux_cond_11_pad;
  wire  mux_cond_12_shl;
  wire [19:0] mux_cond_12_pad;
  wire [13:0] mux_cond_13_shl;
  wire [19:0] mux_cond_13_pad;
  wire [8:0] mux_cond_14_shl;
  wire [19:0] mux_cond_14_pad;
  wire  mux_cond_15_shl;
  wire [19:0] mux_cond_15_pad;
  wire [9:0] mux_cond_16_shl;
  wire [19:0] mux_cond_16_pad;
  wire [13:0] mux_cond_17_shl;
  wire [19:0] mux_cond_17_pad;
  wire [18:0] mux_cond_18_shl;
  wire [19:0] mux_cond_18_pad;
  wire [3:0] mux_cond_19_shl;
  wire [19:0] mux_cond_19_pad;
  wire  mux_cond_20_shl;
  wire [19:0] mux_cond_20_pad;
  wire [10:0] mux_cond_21_shl;
  wire [19:0] mux_cond_21_pad;
  wire [3:0] mux_cond_22_shl;
  wire [19:0] mux_cond_22_pad;
  wire [2:0] mux_cond_23_shl;
  wire [19:0] mux_cond_23_pad;
  wire [7:0] mux_cond_24_shl;
  wire [19:0] mux_cond_24_pad;
  wire [17:0] mux_cond_25_shl;
  wire [19:0] mux_cond_25_pad;
  wire [5:0] mux_cond_26_shl;
  wire [19:0] mux_cond_26_pad;
  wire [6:0] mux_cond_27_shl;
  wire [19:0] mux_cond_27_pad;
  wire [19:0] mux_cond_28_shl;
  wire [19:0] mux_cond_28_pad;
  wire [16:0] mux_cond_29_shl;
  wire [19:0] mux_cond_29_pad;
  wire [18:0] mux_cond_30_shl;
  wire [19:0] mux_cond_30_pad;
  wire  mux_cond_31_shl;
  wire [19:0] mux_cond_31_pad;
  wire [2:0] mux_cond_32_shl;
  wire [19:0] mux_cond_32_pad;
  wire [11:0] mux_cond_33_shl;
  wire [19:0] mux_cond_33_pad;
  wire [18:0] mux_cond_34_shl;
  wire [19:0] mux_cond_34_pad;
  wire [9:0] mux_cond_35_shl;
  wire [19:0] mux_cond_35_pad;
  wire [1:0] mux_cond_36_shl;
  wire [19:0] mux_cond_36_pad;
  wire [1:0] mux_cond_37_shl;
  wire [19:0] mux_cond_37_pad;
  wire [3:0] mux_cond_38_shl;
  wire [19:0] mux_cond_38_pad;
  wire  mux_cond_39_shl;
  wire [19:0] mux_cond_39_pad;
  wire [15:0] mux_cond_40_shl;
  wire [19:0] mux_cond_40_pad;
  wire [6:0] mux_cond_41_shl;
  wire [19:0] mux_cond_41_pad;
  wire [19:0] mux_cond_42_shl;
  wire [19:0] mux_cond_42_pad;
  wire [19:0] mux_cond_43_shl;
  wire [19:0] mux_cond_43_pad;
  wire [13:0] mux_cond_44_shl;
  wire [19:0] mux_cond_44_pad;
  wire [1:0] mux_cond_45_shl;
  wire [19:0] mux_cond_45_pad;
  wire [8:0] mux_cond_46_shl;
  wire [19:0] mux_cond_46_pad;
  wire [17:0] mux_cond_47_shl;
  wire [19:0] mux_cond_47_pad;
  wire [11:0] mux_cond_48_shl;
  wire [19:0] mux_cond_48_pad;
  wire [3:0] mux_cond_49_shl;
  wire [19:0] mux_cond_49_pad;
  wire [11:0] mux_cond_50_shl;
  wire [19:0] mux_cond_50_pad;
  wire [14:0] mux_cond_51_shl;
  wire [19:0] mux_cond_51_pad;
  wire [5:0] mux_cond_52_shl;
  wire [19:0] mux_cond_52_pad;
  wire [3:0] mux_cond_53_shl;
  wire [19:0] mux_cond_53_pad;
  wire [18:0] mux_cond_54_shl;
  wire [19:0] mux_cond_54_pad;
  wire [9:0] mux_cond_55_shl;
  wire [19:0] mux_cond_55_pad;
  wire [15:0] mux_cond_56_shl;
  wire [19:0] mux_cond_56_pad;
  wire [17:0] mux_cond_57_shl;
  wire [19:0] mux_cond_57_pad;
  wire [13:0] mux_cond_58_shl;
  wire [19:0] mux_cond_58_pad;
  wire [12:0] mux_cond_59_shl;
  wire [19:0] mux_cond_59_pad;
  wire [14:0] mux_cond_60_shl;
  wire [19:0] mux_cond_60_pad;
  wire [9:0] mux_cond_61_shl;
  wire [19:0] mux_cond_61_pad;
  wire [4:0] mux_cond_62_shl;
  wire [19:0] mux_cond_62_pad;
  wire [6:0] mux_cond_63_shl;
  wire [19:0] mux_cond_63_pad;
  wire [5:0] mux_cond_64_shl;
  wire [19:0] mux_cond_64_pad;
  wire [9:0] mux_cond_65_shl;
  wire [19:0] mux_cond_65_pad;
  wire  mux_cond_66_shl;
  wire [19:0] mux_cond_66_pad;
  wire [13:0] mux_cond_67_shl;
  wire [19:0] mux_cond_67_pad;
  wire [19:0] mux_cond_68_shl;
  wire [19:0] mux_cond_68_pad;
  wire [8:0] mux_cond_69_shl;
  wire [19:0] mux_cond_69_pad;
  wire [7:0] mux_cond_70_shl;
  wire [19:0] mux_cond_70_pad;
  wire [8:0] mux_cond_71_shl;
  wire [19:0] mux_cond_71_pad;
  wire [3:0] mux_cond_72_shl;
  wire [19:0] mux_cond_72_pad;
  wire [6:0] mux_cond_73_shl;
  wire [19:0] mux_cond_73_pad;
  wire [18:0] mux_cond_74_shl;
  wire [19:0] mux_cond_74_pad;
  wire [18:0] mux_cond_75_shl;
  wire [19:0] mux_cond_75_pad;
  wire [6:0] mux_cond_76_shl;
  wire [19:0] mux_cond_76_pad;
  wire [5:0] mux_cond_77_shl;
  wire [19:0] mux_cond_77_pad;
  wire [14:0] mux_cond_78_shl;
  wire [19:0] mux_cond_78_pad;
  wire [9:0] mux_cond_79_shl;
  wire [19:0] mux_cond_79_pad;
  wire [8:0] mux_cond_80_shl;
  wire [19:0] mux_cond_80_pad;
  wire [10:0] mux_cond_81_shl;
  wire [19:0] mux_cond_81_pad;
  wire [2:0] mux_cond_82_shl;
  wire [19:0] mux_cond_82_pad;
  wire [15:0] mux_cond_83_shl;
  wire [19:0] mux_cond_83_pad;
  wire  mux_cond_84_shl;
  wire [19:0] mux_cond_84_pad;
  wire [1:0] mux_cond_85_shl;
  wire [19:0] mux_cond_85_pad;
  wire [17:0] mux_cond_86_shl;
  wire [19:0] mux_cond_86_pad;
  wire [15:0] mux_cond_87_shl;
  wire [19:0] mux_cond_87_pad;
  wire [14:0] mux_cond_88_shl;
  wire [19:0] mux_cond_88_pad;
  wire [15:0] mux_cond_89_shl;
  wire [19:0] mux_cond_89_pad;
  wire  mux_cond_90_shl;
  wire [19:0] mux_cond_90_pad;
  wire [5:0] mux_cond_91_shl;
  wire [19:0] mux_cond_91_pad;
  wire [19:0] mux_cond_92_shl;
  wire [19:0] mux_cond_92_pad;
  wire [1:0] mux_cond_93_shl;
  wire [19:0] mux_cond_93_pad;
  wire [11:0] mux_cond_94_shl;
  wire [19:0] mux_cond_94_pad;
  wire [8:0] mux_cond_95_shl;
  wire [19:0] mux_cond_95_pad;
  wire [16:0] mux_cond_96_shl;
  wire [19:0] mux_cond_96_pad;
  wire [14:0] mux_cond_97_shl;
  wire [19:0] mux_cond_97_pad;
  wire [19:0] MulDiv_xor64;
  wire [19:0] MulDiv_xor31;
  wire [19:0] MulDiv_xor66;
  wire [19:0] MulDiv_xor32;
  wire [19:0] MulDiv_xor15;
  wire [19:0] MulDiv_xor68;
  wire [19:0] MulDiv_xor33;
  wire [19:0] MulDiv_xor70;
  wire [19:0] MulDiv_xor34;
  wire [19:0] MulDiv_xor16;
  wire [19:0] MulDiv_xor7;
  wire [19:0] MulDiv_xor72;
  wire [19:0] MulDiv_xor35;
  wire [19:0] MulDiv_xor74;
  wire [19:0] MulDiv_xor36;
  wire [19:0] MulDiv_xor17;
  wire [19:0] MulDiv_xor76;
  wire [19:0] MulDiv_xor37;
  wire [19:0] MulDiv_xor77;
  wire [19:0] MulDiv_xor78;
  wire [19:0] MulDiv_xor38;
  wire [19:0] MulDiv_xor18;
  wire [19:0] MulDiv_xor8;
  wire [19:0] MulDiv_xor3;
  wire [19:0] MulDiv_xor80;
  wire [19:0] MulDiv_xor39;
  wire [19:0] MulDiv_xor82;
  wire [19:0] MulDiv_xor40;
  wire [19:0] MulDiv_xor19;
  wire [19:0] MulDiv_xor84;
  wire [19:0] MulDiv_xor41;
  wire [19:0] MulDiv_xor85;
  wire [19:0] MulDiv_xor86;
  wire [19:0] MulDiv_xor42;
  wire [19:0] MulDiv_xor20;
  wire [19:0] MulDiv_xor9;
  wire [19:0] MulDiv_xor88;
  wire [19:0] MulDiv_xor43;
  wire [19:0] MulDiv_xor90;
  wire [19:0] MulDiv_xor44;
  wire [19:0] MulDiv_xor21;
  wire [19:0] MulDiv_xor92;
  wire [19:0] MulDiv_xor45;
  wire [19:0] MulDiv_xor93;
  wire [19:0] MulDiv_xor94;
  wire [19:0] MulDiv_xor46;
  wire [19:0] MulDiv_xor22;
  wire [19:0] MulDiv_xor10;
  wire [19:0] MulDiv_xor4;
  wire [19:0] MulDiv_xor1;
  wire [19:0] MulDiv_xor96;
  wire [19:0] MulDiv_xor47;
  wire [19:0] MulDiv_xor98;
  wire [19:0] MulDiv_xor48;
  wire [19:0] MulDiv_xor23;
  wire [19:0] MulDiv_xor100;
  wire [19:0] MulDiv_xor49;
  wire [19:0] MulDiv_xor101;
  wire [19:0] MulDiv_xor102;
  wire [19:0] MulDiv_xor50;
  wire [19:0] MulDiv_xor24;
  wire [19:0] MulDiv_xor11;
  wire [19:0] MulDiv_xor104;
  wire [19:0] MulDiv_xor51;
  wire [19:0] MulDiv_xor106;
  wire [19:0] MulDiv_xor52;
  wire [19:0] MulDiv_xor25;
  wire [19:0] MulDiv_xor108;
  wire [19:0] MulDiv_xor53;
  wire [19:0] MulDiv_xor109;
  wire [19:0] MulDiv_xor110;
  wire [19:0] MulDiv_xor54;
  wire [19:0] MulDiv_xor26;
  wire [19:0] MulDiv_xor12;
  wire [19:0] MulDiv_xor5;
  wire [19:0] MulDiv_xor112;
  wire [19:0] MulDiv_xor55;
  wire [19:0] MulDiv_xor114;
  wire [19:0] MulDiv_xor56;
  wire [19:0] MulDiv_xor27;
  wire [19:0] MulDiv_xor116;
  wire [19:0] MulDiv_xor57;
  wire [19:0] MulDiv_xor117;
  wire [19:0] MulDiv_xor118;
  wire [19:0] MulDiv_xor58;
  wire [19:0] MulDiv_xor28;
  wire [19:0] MulDiv_xor13;
  wire [19:0] MulDiv_xor120;
  wire [19:0] MulDiv_xor59;
  wire [19:0] MulDiv_xor122;
  wire [19:0] MulDiv_xor60;
  wire [19:0] MulDiv_xor29;
  wire [19:0] MulDiv_xor124;
  wire [19:0] MulDiv_xor61;
  wire [19:0] MulDiv_xor125;
  wire [19:0] MulDiv_xor126;
  wire [19:0] MulDiv_xor62;
  wire [19:0] MulDiv_xor30;
  wire [19:0] MulDiv_xor14;
  wire [19:0] MulDiv_xor6;
  wire [19:0] MulDiv_xor2;
  wire [19:0] MulDiv_xor0;
  assign _T_22 = io_req_bits_fn & 4'h4; // @[Decode.scala 14:65]
  assign cmdMul = _T_22 == 4'h0; // @[Decode.scala 14:121]
  assign _T_25 = io_req_bits_fn & 4'h5; // @[Decode.scala 14:65]
  assign _T_26 = _T_25 == 4'h1; // @[Decode.scala 14:121]
  assign _T_27 = io_req_bits_fn & 4'h2; // @[Decode.scala 14:65]
  assign _T_28 = _T_27 == 4'h2; // @[Decode.scala 14:121]
  assign cmdHi = _T_26 | _T_28; // @[Decode.scala 15:30]
  assign _T_31 = io_req_bits_fn & 4'h6; // @[Decode.scala 14:65]
  assign _T_32 = _T_31 == 4'h0; // @[Decode.scala 14:121]
  assign _T_33 = io_req_bits_fn & 4'h1; // @[Decode.scala 14:65]
  assign _T_34 = _T_33 == 4'h0; // @[Decode.scala 14:121]
  assign lhsSigned = _T_32 | _T_34; // @[Decode.scala 15:30]
  assign _T_38 = _T_25 == 4'h4; // @[Decode.scala 14:121]
  assign rhsSigned = _T_32 | _T_38; // @[Decode.scala 15:30]
  assign _T_45 = io_req_bits_dw ? io_req_bits_in1[63] : io_req_bits_in1[31]; // @[Multiplier.scala 81:29]
  assign lhs_sign = lhsSigned & _T_45; // @[Multiplier.scala 81:23]
  assign _T_47 = lhs_sign ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  assign _T_49 = io_req_bits_dw ? io_req_bits_in1[63:32] : _T_47; // @[Multiplier.scala 82:17]
  assign lhs_in = {_T_49,io_req_bits_in1[31:0]}; // @[Cat.scala 30:58]
  assign _T_55 = io_req_bits_dw ? io_req_bits_in2[63] : io_req_bits_in2[31]; // @[Multiplier.scala 81:29]
  assign rhs_sign = rhsSigned & _T_55; // @[Multiplier.scala 81:23]
  assign _T_57 = rhs_sign ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  assign _T_59 = io_req_bits_dw ? io_req_bits_in2[63:32] : _T_57; // @[Multiplier.scala 82:17]
  assign subtractor = remainder[128:64] - divisor; // @[Multiplier.scala 88:37]
  assign result = resHi ? remainder[128:65] : remainder[63:0]; // @[Multiplier.scala 89:19]
  assign negated_remainder = 64'h0 - result; // @[Multiplier.scala 90:27]
  assign _T_68 = state == 3'h1; // @[Multiplier.scala 92:39]
  assign _T_71 = state == 3'h5; // @[Multiplier.scala 101:39]
  assign _T_72 = state == 3'h2; // @[Multiplier.scala 106:39]
  assign _T_75 = {remainder[129:65],remainder[63:0]}; // @[Cat.scala 30:58]
  assign _T_79 = _T_75[128:64]; // @[Multiplier.scala 110:37]
  assign _T_83 = {remainder[64],_T_75[7:0]}; // @[Multiplier.scala 112:60]
  assign _GEN_37 = {{56{_T_83[8]}},_T_83}; // @[Multiplier.scala 112:67]
  assign _T_84 = $signed(_GEN_37) * $signed(divisor); // @[Multiplier.scala 112:67]
  assign _GEN_38 = {{9{_T_79[64]}},_T_79}; // @[Multiplier.scala 112:76]
  assign _T_89 = $signed(_T_84) + $signed(_GEN_38); // @[Cat.scala 30:58]
  assign _T_90 = {_T_89,_T_75[63:8]}; // @[Cat.scala 30:58]
  assign _T_91 = count == 7'h6; // @[Multiplier.scala 114:32]
  assign _T_92 = _T_91 & neg_out; // @[Multiplier.scala 114:57]
  assign _T_93 = count * 7'h8; // @[Multiplier.scala 116:56]
  assign _T_95 = -65'sh10000000000000000 >>> _T_93[5:0]; // @[Multiplier.scala 116:46]
  assign _T_97 = count != 7'h7; // @[Multiplier.scala 117:47]
  assign _T_99 = count != 7'h0; // @[Multiplier.scala 117:81]
  assign _T_100 = _T_97 & _T_99; // @[Multiplier.scala 117:72]
  assign _T_102 = _T_100 & ~isHi; // @[Multiplier.scala 117:87]
  assign _T_104 = _T_75[63:0] & ~_T_95[63:0]; // @[Multiplier.scala 118:24]
  assign _T_105 = _T_104 == 64'h0; // @[Multiplier.scala 118:37]
  assign _T_106 = _T_102 & _T_105; // @[Multiplier.scala 118:13]
  assign _T_110 = 11'h40 - _T_93; // @[Multiplier.scala 119:36]
  assign _T_112 = _T_75 >> _T_110[5:0]; // @[Multiplier.scala 119:27]
  assign _T_114 = _T_106 ? {{1'd0}, _T_112} : _T_90; // @[Multiplier.scala 120:55]
  assign _T_116 = {_T_90[128:64],_T_114[63:0]}; // @[Cat.scala 30:58]
  assign _T_120 = {_T_116[128:64],_T_92,_T_116[63:0]}; // @[Cat.scala 30:58]
  assign _T_122 = count + 7'h1; // @[Multiplier.scala 123:20]
  assign _T_123 = count == 7'h7; // @[Multiplier.scala 124:25]
  assign _T_124 = _T_106 | _T_123; // @[Multiplier.scala 124:16]
  assign _T_125 = state == 3'h3; // @[Multiplier.scala 129:39]
  assign _T_129 = subtractor[64] ? remainder[127:64] : subtractor[63:0]; // @[Multiplier.scala 134:14]
  assign _T_133 = {_T_129,remainder[63:0],~subtractor[64]}; // @[Cat.scala 30:58]
  assign _T_134 = count == 7'h40; // @[Multiplier.scala 138:17]
  assign _T_138 = count == 7'h0; // @[Multiplier.scala 146:24]
  assign _T_141 = _T_138 & ~subtractor[64]; // @[Multiplier.scala 146:30]
  assign _T_146 = divisor[63:32] != 32'h0; // @[CircuitMath.scala 37:22]
  assign _T_149 = divisor[63:48] != 16'h0; // @[CircuitMath.scala 37:22]
  assign _T_152 = divisor[63:56] != 8'h0; // @[CircuitMath.scala 37:22]
  assign _T_155 = divisor[63:60] != 4'h0; // @[CircuitMath.scala 37:22]
  assign _T_159 = divisor[62] ? 2'h2 : {{1'd0}, divisor[61]}; // @[CircuitMath.scala 32:10]
  assign _T_160 = divisor[63] ? 2'h3 : _T_159; // @[CircuitMath.scala 32:10]
  assign _T_164 = divisor[58] ? 2'h2 : {{1'd0}, divisor[57]}; // @[CircuitMath.scala 32:10]
  assign _T_165 = divisor[59] ? 2'h3 : _T_164; // @[CircuitMath.scala 32:10]
  assign _T_166 = _T_155 ? _T_160 : _T_165; // @[CircuitMath.scala 38:21]
  assign _T_167 = {_T_155,_T_166}; // @[Cat.scala 30:58]
  assign _T_170 = divisor[55:52] != 4'h0; // @[CircuitMath.scala 37:22]
  assign _T_174 = divisor[54] ? 2'h2 : {{1'd0}, divisor[53]}; // @[CircuitMath.scala 32:10]
  assign _T_175 = divisor[55] ? 2'h3 : _T_174; // @[CircuitMath.scala 32:10]
  assign _T_179 = divisor[50] ? 2'h2 : {{1'd0}, divisor[49]}; // @[CircuitMath.scala 32:10]
  assign _T_180 = divisor[51] ? 2'h3 : _T_179; // @[CircuitMath.scala 32:10]
  assign _T_181 = _T_170 ? _T_175 : _T_180; // @[CircuitMath.scala 38:21]
  assign _T_182 = {_T_170,_T_181}; // @[Cat.scala 30:58]
  assign _T_183 = _T_152 ? _T_167 : _T_182; // @[CircuitMath.scala 38:21]
  assign _T_184 = {_T_152,_T_183}; // @[Cat.scala 30:58]
  assign _T_187 = divisor[47:40] != 8'h0; // @[CircuitMath.scala 37:22]
  assign _T_190 = divisor[47:44] != 4'h0; // @[CircuitMath.scala 37:22]
  assign _T_194 = divisor[46] ? 2'h2 : {{1'd0}, divisor[45]}; // @[CircuitMath.scala 32:10]
  assign _T_195 = divisor[47] ? 2'h3 : _T_194; // @[CircuitMath.scala 32:10]
  assign _T_199 = divisor[42] ? 2'h2 : {{1'd0}, divisor[41]}; // @[CircuitMath.scala 32:10]
  assign _T_200 = divisor[43] ? 2'h3 : _T_199; // @[CircuitMath.scala 32:10]
  assign _T_201 = _T_190 ? _T_195 : _T_200; // @[CircuitMath.scala 38:21]
  assign _T_202 = {_T_190,_T_201}; // @[Cat.scala 30:58]
  assign _T_205 = divisor[39:36] != 4'h0; // @[CircuitMath.scala 37:22]
  assign _T_209 = divisor[38] ? 2'h2 : {{1'd0}, divisor[37]}; // @[CircuitMath.scala 32:10]
  assign _T_210 = divisor[39] ? 2'h3 : _T_209; // @[CircuitMath.scala 32:10]
  assign _T_214 = divisor[34] ? 2'h2 : {{1'd0}, divisor[33]}; // @[CircuitMath.scala 32:10]
  assign _T_215 = divisor[35] ? 2'h3 : _T_214; // @[CircuitMath.scala 32:10]
  assign _T_216 = _T_205 ? _T_210 : _T_215; // @[CircuitMath.scala 38:21]
  assign _T_217 = {_T_205,_T_216}; // @[Cat.scala 30:58]
  assign _T_218 = _T_187 ? _T_202 : _T_217; // @[CircuitMath.scala 38:21]
  assign _T_219 = {_T_187,_T_218}; // @[Cat.scala 30:58]
  assign _T_220 = _T_149 ? _T_184 : _T_219; // @[CircuitMath.scala 38:21]
  assign _T_221 = {_T_149,_T_220}; // @[Cat.scala 30:58]
  assign _T_224 = divisor[31:16] != 16'h0; // @[CircuitMath.scala 37:22]
  assign _T_227 = divisor[31:24] != 8'h0; // @[CircuitMath.scala 37:22]
  assign _T_230 = divisor[31:28] != 4'h0; // @[CircuitMath.scala 37:22]
  assign _T_234 = divisor[30] ? 2'h2 : {{1'd0}, divisor[29]}; // @[CircuitMath.scala 32:10]
  assign _T_235 = divisor[31] ? 2'h3 : _T_234; // @[CircuitMath.scala 32:10]
  assign _T_239 = divisor[26] ? 2'h2 : {{1'd0}, divisor[25]}; // @[CircuitMath.scala 32:10]
  assign _T_240 = divisor[27] ? 2'h3 : _T_239; // @[CircuitMath.scala 32:10]
  assign _T_241 = _T_230 ? _T_235 : _T_240; // @[CircuitMath.scala 38:21]
  assign _T_242 = {_T_230,_T_241}; // @[Cat.scala 30:58]
  assign _T_245 = divisor[23:20] != 4'h0; // @[CircuitMath.scala 37:22]
  assign _T_249 = divisor[22] ? 2'h2 : {{1'd0}, divisor[21]}; // @[CircuitMath.scala 32:10]
  assign _T_250 = divisor[23] ? 2'h3 : _T_249; // @[CircuitMath.scala 32:10]
  assign _T_254 = divisor[18] ? 2'h2 : {{1'd0}, divisor[17]}; // @[CircuitMath.scala 32:10]
  assign _T_255 = divisor[19] ? 2'h3 : _T_254; // @[CircuitMath.scala 32:10]
  assign _T_256 = _T_245 ? _T_250 : _T_255; // @[CircuitMath.scala 38:21]
  assign _T_257 = {_T_245,_T_256}; // @[Cat.scala 30:58]
  assign _T_258 = _T_227 ? _T_242 : _T_257; // @[CircuitMath.scala 38:21]
  assign _T_259 = {_T_227,_T_258}; // @[Cat.scala 30:58]
  assign _T_262 = divisor[15:8] != 8'h0; // @[CircuitMath.scala 37:22]
  assign _T_265 = divisor[15:12] != 4'h0; // @[CircuitMath.scala 37:22]
  assign _T_269 = divisor[14] ? 2'h2 : {{1'd0}, divisor[13]}; // @[CircuitMath.scala 32:10]
  assign _T_270 = divisor[15] ? 2'h3 : _T_269; // @[CircuitMath.scala 32:10]
  assign _T_274 = divisor[10] ? 2'h2 : {{1'd0}, divisor[9]}; // @[CircuitMath.scala 32:10]
  assign _T_275 = divisor[11] ? 2'h3 : _T_274; // @[CircuitMath.scala 32:10]
  assign _T_276 = _T_265 ? _T_270 : _T_275; // @[CircuitMath.scala 38:21]
  assign _T_277 = {_T_265,_T_276}; // @[Cat.scala 30:58]
  assign _T_280 = divisor[7:4] != 4'h0; // @[CircuitMath.scala 37:22]
  assign _T_284 = divisor[6] ? 2'h2 : {{1'd0}, divisor[5]}; // @[CircuitMath.scala 32:10]
  assign _T_285 = divisor[7] ? 2'h3 : _T_284; // @[CircuitMath.scala 32:10]
  assign _T_289 = divisor[2] ? 2'h2 : {{1'd0}, divisor[1]}; // @[CircuitMath.scala 32:10]
  assign _T_290 = divisor[3] ? 2'h3 : _T_289; // @[CircuitMath.scala 32:10]
  assign _T_291 = _T_280 ? _T_285 : _T_290; // @[CircuitMath.scala 38:21]
  assign _T_292 = {_T_280,_T_291}; // @[Cat.scala 30:58]
  assign _T_293 = _T_262 ? _T_277 : _T_292; // @[CircuitMath.scala 38:21]
  assign _T_294 = {_T_262,_T_293}; // @[Cat.scala 30:58]
  assign _T_295 = _T_224 ? _T_259 : _T_294; // @[CircuitMath.scala 38:21]
  assign _T_296 = {_T_224,_T_295}; // @[Cat.scala 30:58]
  assign _T_297 = _T_146 ? _T_221 : _T_296; // @[CircuitMath.scala 38:21]
  assign _T_298 = {_T_146,_T_297}; // @[Cat.scala 30:58]
  assign _T_303 = remainder[63:32] != 32'h0; // @[CircuitMath.scala 37:22]
  assign _T_306 = remainder[63:48] != 16'h0; // @[CircuitMath.scala 37:22]
  assign _T_309 = remainder[63:56] != 8'h0; // @[CircuitMath.scala 37:22]
  assign _T_312 = remainder[63:60] != 4'h0; // @[CircuitMath.scala 37:22]
  assign _T_316 = remainder[62] ? 2'h2 : {{1'd0}, remainder[61]}; // @[CircuitMath.scala 32:10]
  assign _T_317 = remainder[63] ? 2'h3 : _T_316; // @[CircuitMath.scala 32:10]
  assign _T_321 = remainder[58] ? 2'h2 : {{1'd0}, remainder[57]}; // @[CircuitMath.scala 32:10]
  assign _T_322 = remainder[59] ? 2'h3 : _T_321; // @[CircuitMath.scala 32:10]
  assign _T_323 = _T_312 ? _T_317 : _T_322; // @[CircuitMath.scala 38:21]
  assign _T_324 = {_T_312,_T_323}; // @[Cat.scala 30:58]
  assign _T_327 = remainder[55:52] != 4'h0; // @[CircuitMath.scala 37:22]
  assign _T_331 = remainder[54] ? 2'h2 : {{1'd0}, remainder[53]}; // @[CircuitMath.scala 32:10]
  assign _T_332 = remainder[55] ? 2'h3 : _T_331; // @[CircuitMath.scala 32:10]
  assign _T_336 = remainder[50] ? 2'h2 : {{1'd0}, remainder[49]}; // @[CircuitMath.scala 32:10]
  assign _T_337 = remainder[51] ? 2'h3 : _T_336; // @[CircuitMath.scala 32:10]
  assign _T_338 = _T_327 ? _T_332 : _T_337; // @[CircuitMath.scala 38:21]
  assign _T_339 = {_T_327,_T_338}; // @[Cat.scala 30:58]
  assign _T_340 = _T_309 ? _T_324 : _T_339; // @[CircuitMath.scala 38:21]
  assign _T_341 = {_T_309,_T_340}; // @[Cat.scala 30:58]
  assign _T_344 = remainder[47:40] != 8'h0; // @[CircuitMath.scala 37:22]
  assign _T_347 = remainder[47:44] != 4'h0; // @[CircuitMath.scala 37:22]
  assign _T_351 = remainder[46] ? 2'h2 : {{1'd0}, remainder[45]}; // @[CircuitMath.scala 32:10]
  assign _T_352 = remainder[47] ? 2'h3 : _T_351; // @[CircuitMath.scala 32:10]
  assign _T_356 = remainder[42] ? 2'h2 : {{1'd0}, remainder[41]}; // @[CircuitMath.scala 32:10]
  assign _T_357 = remainder[43] ? 2'h3 : _T_356; // @[CircuitMath.scala 32:10]
  assign _T_358 = _T_347 ? _T_352 : _T_357; // @[CircuitMath.scala 38:21]
  assign _T_359 = {_T_347,_T_358}; // @[Cat.scala 30:58]
  assign _T_362 = remainder[39:36] != 4'h0; // @[CircuitMath.scala 37:22]
  assign _T_366 = remainder[38] ? 2'h2 : {{1'd0}, remainder[37]}; // @[CircuitMath.scala 32:10]
  assign _T_367 = remainder[39] ? 2'h3 : _T_366; // @[CircuitMath.scala 32:10]
  assign _T_371 = remainder[34] ? 2'h2 : {{1'd0}, remainder[33]}; // @[CircuitMath.scala 32:10]
  assign _T_372 = remainder[35] ? 2'h3 : _T_371; // @[CircuitMath.scala 32:10]
  assign _T_373 = _T_362 ? _T_367 : _T_372; // @[CircuitMath.scala 38:21]
  assign _T_374 = {_T_362,_T_373}; // @[Cat.scala 30:58]
  assign _T_375 = _T_344 ? _T_359 : _T_374; // @[CircuitMath.scala 38:21]
  assign _T_376 = {_T_344,_T_375}; // @[Cat.scala 30:58]
  assign _T_377 = _T_306 ? _T_341 : _T_376; // @[CircuitMath.scala 38:21]
  assign _T_378 = {_T_306,_T_377}; // @[Cat.scala 30:58]
  assign _T_381 = remainder[31:16] != 16'h0; // @[CircuitMath.scala 37:22]
  assign _T_384 = remainder[31:24] != 8'h0; // @[CircuitMath.scala 37:22]
  assign _T_387 = remainder[31:28] != 4'h0; // @[CircuitMath.scala 37:22]
  assign _T_391 = remainder[30] ? 2'h2 : {{1'd0}, remainder[29]}; // @[CircuitMath.scala 32:10]
  assign _T_392 = remainder[31] ? 2'h3 : _T_391; // @[CircuitMath.scala 32:10]
  assign _T_396 = remainder[26] ? 2'h2 : {{1'd0}, remainder[25]}; // @[CircuitMath.scala 32:10]
  assign _T_397 = remainder[27] ? 2'h3 : _T_396; // @[CircuitMath.scala 32:10]
  assign _T_398 = _T_387 ? _T_392 : _T_397; // @[CircuitMath.scala 38:21]
  assign _T_399 = {_T_387,_T_398}; // @[Cat.scala 30:58]
  assign _T_402 = remainder[23:20] != 4'h0; // @[CircuitMath.scala 37:22]
  assign _T_406 = remainder[22] ? 2'h2 : {{1'd0}, remainder[21]}; // @[CircuitMath.scala 32:10]
  assign _T_407 = remainder[23] ? 2'h3 : _T_406; // @[CircuitMath.scala 32:10]
  assign _T_411 = remainder[18] ? 2'h2 : {{1'd0}, remainder[17]}; // @[CircuitMath.scala 32:10]
  assign _T_412 = remainder[19] ? 2'h3 : _T_411; // @[CircuitMath.scala 32:10]
  assign _T_413 = _T_402 ? _T_407 : _T_412; // @[CircuitMath.scala 38:21]
  assign _T_414 = {_T_402,_T_413}; // @[Cat.scala 30:58]
  assign _T_415 = _T_384 ? _T_399 : _T_414; // @[CircuitMath.scala 38:21]
  assign _T_416 = {_T_384,_T_415}; // @[Cat.scala 30:58]
  assign _T_419 = remainder[15:8] != 8'h0; // @[CircuitMath.scala 37:22]
  assign _T_422 = remainder[15:12] != 4'h0; // @[CircuitMath.scala 37:22]
  assign _T_426 = remainder[14] ? 2'h2 : {{1'd0}, remainder[13]}; // @[CircuitMath.scala 32:10]
  assign _T_427 = remainder[15] ? 2'h3 : _T_426; // @[CircuitMath.scala 32:10]
  assign _T_431 = remainder[10] ? 2'h2 : {{1'd0}, remainder[9]}; // @[CircuitMath.scala 32:10]
  assign _T_432 = remainder[11] ? 2'h3 : _T_431; // @[CircuitMath.scala 32:10]
  assign _T_433 = _T_422 ? _T_427 : _T_432; // @[CircuitMath.scala 38:21]
  assign _T_434 = {_T_422,_T_433}; // @[Cat.scala 30:58]
  assign _T_437 = remainder[7:4] != 4'h0; // @[CircuitMath.scala 37:22]
  assign _T_441 = remainder[6] ? 2'h2 : {{1'd0}, remainder[5]}; // @[CircuitMath.scala 32:10]
  assign _T_442 = remainder[7] ? 2'h3 : _T_441; // @[CircuitMath.scala 32:10]
  assign _T_446 = remainder[2] ? 2'h2 : {{1'd0}, remainder[1]}; // @[CircuitMath.scala 32:10]
  assign _T_447 = remainder[3] ? 2'h3 : _T_446; // @[CircuitMath.scala 32:10]
  assign _T_448 = _T_437 ? _T_442 : _T_447; // @[CircuitMath.scala 38:21]
  assign _T_449 = {_T_437,_T_448}; // @[Cat.scala 30:58]
  assign _T_450 = _T_419 ? _T_434 : _T_449; // @[CircuitMath.scala 38:21]
  assign _T_451 = {_T_419,_T_450}; // @[Cat.scala 30:58]
  assign _T_452 = _T_381 ? _T_416 : _T_451; // @[CircuitMath.scala 38:21]
  assign _T_453 = {_T_381,_T_452}; // @[Cat.scala 30:58]
  assign _T_454 = _T_303 ? _T_378 : _T_453; // @[CircuitMath.scala 38:21]
  assign _T_455 = {_T_303,_T_454}; // @[Cat.scala 30:58]
  assign _T_460 = _T_455 - _T_298; // @[Multiplier.scala 152:35]
  assign _T_464 = _T_138 & ~_T_141; // @[Multiplier.scala 153:30]
  assign _T_465 = ~_T_460 >= 6'h1; // @[Multiplier.scala 153:52]
  assign _T_466 = _T_464 & _T_465; // @[Multiplier.scala 153:41]
  assign _GEN_39 = {{63'd0}, remainder[63:0]}; // @[Multiplier.scala 155:39]
  assign _T_468 = _GEN_39 << ~_T_460; // @[Multiplier.scala 155:39]
  assign _GEN_16 = _T_466 ? {{2'd0}, _T_468} : _T_133; // @[Multiplier.scala 154:19]
  assign _T_471 = _T_141 & ~isHi; // @[Multiplier.scala 159:18]
  assign _T_472 = io_resp_ready & io_resp_valid; // @[Decoupled.scala 37:37]
  assign _T_473 = _T_472 | io_kill; // @[Multiplier.scala 161:24]
  assign _T_474 = io_req_ready & io_req_valid; // @[Decoupled.scala 37:37]
  assign _T_475 = lhs_sign | rhs_sign; // @[Multiplier.scala 165:46]
  assign _T_480 = cmdMul & ~io_req_bits_dw; // @[Multiplier.scala 168:46]
  assign _T_481 = _T_480 ? 3'h4 : 3'h0; // @[Multiplier.scala 168:38]
  assign _T_482 = lhs_sign != rhs_sign; // @[Multiplier.scala 169:46]
  assign _T_484 = {rhs_sign,_T_59,io_req_bits_in2[31:0]}; // @[Cat.scala 30:58]
  assign _T_486 = state & 3'h1; // @[Multiplier.scala 175:23]
  assign outMul = _T_486 == 3'h0; // @[Multiplier.scala 175:52]
  assign _T_492 = ~req_dw & outMul; // @[Multiplier.scala 176:52]
  assign loOut = _T_492 ? result[63:32] : result[31:0]; // @[Multiplier.scala 176:18]
  assign _T_499 = loOut[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  assign hiOut = req_dw ? result[63:32] : _T_499; // @[Multiplier.scala 177:18]
  assign _T_502 = state == 3'h6; // @[Multiplier.scala 180:27]
  assign _T_503 = state == 3'h7; // @[Multiplier.scala 180:51]
  assign io_req_ready = state == 3'h0; // @[Multiplier.scala 181:16]
  assign io_resp_valid = _T_502 | _T_503; // @[Multiplier.scala 180:17]
  assign io_resp_bits_data = {hiOut,loOut}; // @[Multiplier.scala 179:21]
  assign io_resp_bits_tag = req_tag; // @[Multiplier.scala 178:16]
  assign MulDiv_cov_read_addr = MulDiv_state;
  assign MulDiv_cov_read_data = MulDiv_cov[MulDiv_cov_read_addr]; // @[Coverage map for MulDiv]
  assign MulDiv_cov_write_data = 1'h1;
  assign MulDiv_cov_write_addr = MulDiv_state;
  assign MulDiv_cov_write_mask = 1'h1;
  assign MulDiv_cov_write_en = 1'h1;
  assign mux_cond_0 = _T_347;
  assign mux_cond_1 = _T_205;
  assign mux_cond_2 = remainder[30];
  assign mux_cond_3 = _T_303;
  assign mux_cond_4 = divisor[2];
  assign mux_cond_5 = _T_265;
  assign mux_cond_6 = divisor[38];
  assign mux_cond_7 = _T_419;
  assign mux_cond_8 = divisor[7];
  assign mux_cond_9 = _T_230;
  assign mux_cond_10 = remainder[63];
  assign mux_cond_11 = remainder[6];
  assign mux_cond_12 = loOut[31];
  assign mux_cond_13 = remainder[34];
  assign mux_cond_14 = _T_306;
  assign mux_cond_15 = _T_280;
  assign mux_cond_16 = divisor[62];
  assign mux_cond_17 = remainder[7];
  assign mux_cond_18 = remainder[2];
  assign mux_cond_19 = _T_227;
  assign mux_cond_20 = remainder[31];
  assign mux_cond_21 = remainder[11];
  assign mux_cond_22 = remainder[15];
  assign mux_cond_23 = divisor[42];
  assign mux_cond_24 = divisor[18];
  assign mux_cond_25 = remainder[58];
  assign mux_cond_26 = _T_402;
  assign mux_cond_27 = divisor[59];
  assign mux_cond_28 = remainder[3];
  assign mux_cond_29 = _T_152;
  assign mux_cond_30 = divisor[19];
  assign mux_cond_31 = _T_437;
  assign mux_cond_32 = divisor[35];
  assign mux_cond_33 = divisor[43];
  assign mux_cond_34 = remainder[35];
  assign mux_cond_35 = _T_387;
  assign mux_cond_36 = subtractor[64];
  assign mux_cond_37 = divisor[51];
  assign mux_cond_38 = divisor[58];
  assign mux_cond_39 = remainder[27];
  assign mux_cond_40 = remainder[39];
  assign mux_cond_41 = divisor[47];
  assign mux_cond_42 = _T_422;
  assign mux_cond_43 = divisor[15];
  assign mux_cond_44 = _T_384;
  assign mux_cond_45 = divisor[14];
  assign mux_cond_46 = remainder[23];
  assign mux_cond_47 = divisor[27];
  assign mux_cond_48 = _T_344;
  assign mux_cond_49 = _T_155;
  assign mux_cond_50 = divisor[6];
  assign mux_cond_51 = _T_224;
  assign mux_cond_52 = divisor[63];
  assign mux_cond_53 = remainder[63];
  assign mux_cond_54 = divisor[34];
  assign mux_cond_55 = divisor[46];
  assign mux_cond_56 = _T_245;
  assign mux_cond_57 = divisor[10];
  assign mux_cond_58 = divisor[23];
  assign mux_cond_59 = _T_190;
  assign mux_cond_60 = divisor[3];
  assign mux_cond_61 = remainder[46];
  assign mux_cond_62 = _T_187;
  assign mux_cond_63 = _T_381;
  assign mux_cond_64 = divisor[30];
  assign mux_cond_65 = _T_312;
  assign mux_cond_66 = divisor[11];
  assign mux_cond_67 = divisor[55];
  assign mux_cond_68 = remainder[38];
  assign mux_cond_69 = remainder[43];
  assign mux_cond_70 = remainder[14];
  assign mux_cond_71 = _T_170;
  assign mux_cond_72 = remainder[19];
  assign mux_cond_73 = remainder[62];
  assign mux_cond_74 = divisor[39];
  assign mux_cond_75 = _T_362;
  assign mux_cond_76 = _T_146;
  assign mux_cond_77 = _T_327;
  assign mux_cond_78 = _T_309;
  assign mux_cond_79 = _T_149;
  assign mux_cond_80 = divisor[31];
  assign mux_cond_81 = remainder[47];
  assign mux_cond_82 = remainder[18];
  assign mux_cond_83 = remainder[50];
  assign mux_cond_84 = divisor[22];
  assign mux_cond_85 = remainder[51];
  assign mux_cond_86 = remainder[22];
  assign mux_cond_87 = remainder[55];
  assign mux_cond_88 = remainder[54];
  assign mux_cond_89 = divisor[54];
  assign mux_cond_90 = remainder[26];
  assign mux_cond_91 = _T_262;
  assign mux_cond_92 = remainder[59];
  assign mux_cond_93 = divisor[50];
  assign mux_cond_94 = remainder[42];
  assign mux_cond_95 = remainder[10];
  assign mux_cond_96 = divisor[26];
  assign mux_cond_97 = divisor[63];
  assign resHi_shl = {resHi, 10'h0};
  assign resHi_pad = {9'h0,resHi_shl};
  assign state_shl = {state, 11'h0};
  assign state_pad = {6'h0,state_shl};
  assign req_dw_shl = {req_dw, 5'h0};
  assign req_dw_pad = {14'h0,req_dw_shl};
  assign neg_out_shl = {neg_out, 16'h0};
  assign neg_out_pad = {3'h0,neg_out_shl};
  assign isHi_shl = {isHi, 13'h0};
  assign isHi_pad = {6'h0,isHi_shl};
  assign mux_cond_0_shl = {mux_cond_0, 8'h0};
  assign mux_cond_0_pad = {11'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = mux_cond_1;
  assign mux_cond_1_pad = {19'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 11'h0};
  assign mux_cond_2_pad = {8'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 9'h0};
  assign mux_cond_3_pad = {10'h0,mux_cond_3_shl};
  assign mux_cond_4_shl = {mux_cond_4, 7'h0};
  assign mux_cond_4_pad = {12'h0,mux_cond_4_shl};
  assign mux_cond_5_shl = {mux_cond_5, 5'h0};
  assign mux_cond_5_pad = {14'h0,mux_cond_5_shl};
  assign mux_cond_6_shl = {mux_cond_6, 12'h0};
  assign mux_cond_6_pad = {7'h0,mux_cond_6_shl};
  assign mux_cond_7_shl = {mux_cond_7, 9'h0};
  assign mux_cond_7_pad = {10'h0,mux_cond_7_shl};
  assign mux_cond_8_shl = {mux_cond_8, 2'h0};
  assign mux_cond_8_pad = {17'h0,mux_cond_8_shl};
  assign mux_cond_9_shl = {mux_cond_9, 1'h0};
  assign mux_cond_9_pad = {18'h0,mux_cond_9_shl};
  assign mux_cond_10_shl = {mux_cond_10, 12'h0};
  assign mux_cond_10_pad = {7'h0,mux_cond_10_shl};
  assign mux_cond_11_shl = {mux_cond_11, 8'h0};
  assign mux_cond_11_pad = {11'h0,mux_cond_11_shl};
  assign mux_cond_12_shl = mux_cond_12;
  assign mux_cond_12_pad = {19'h0,mux_cond_12_shl};
  assign mux_cond_13_shl = {mux_cond_13, 13'h0};
  assign mux_cond_13_pad = {6'h0,mux_cond_13_shl};
  assign mux_cond_14_shl = {mux_cond_14, 8'h0};
  assign mux_cond_14_pad = {11'h0,mux_cond_14_shl};
  assign mux_cond_15_shl = mux_cond_15;
  assign mux_cond_15_pad = {19'h0,mux_cond_15_shl};
  assign mux_cond_16_shl = {mux_cond_16, 9'h0};
  assign mux_cond_16_pad = {10'h0,mux_cond_16_shl};
  assign mux_cond_17_shl = {mux_cond_17, 13'h0};
  assign mux_cond_17_pad = {6'h0,mux_cond_17_shl};
  assign mux_cond_18_shl = {mux_cond_18, 18'h0};
  assign mux_cond_18_pad = {1'h0,mux_cond_18_shl};
  assign mux_cond_19_shl = {mux_cond_19, 3'h0};
  assign mux_cond_19_pad = {16'h0,mux_cond_19_shl};
  assign mux_cond_20_shl = mux_cond_20;
  assign mux_cond_20_pad = {19'h0,mux_cond_20_shl};
  assign mux_cond_21_shl = {mux_cond_21, 10'h0};
  assign mux_cond_21_pad = {9'h0,mux_cond_21_shl};
  assign mux_cond_22_shl = {mux_cond_22, 3'h0};
  assign mux_cond_22_pad = {16'h0,mux_cond_22_shl};
  assign mux_cond_23_shl = {mux_cond_23, 2'h0};
  assign mux_cond_23_pad = {17'h0,mux_cond_23_shl};
  assign mux_cond_24_shl = {mux_cond_24, 7'h0};
  assign mux_cond_24_pad = {12'h0,mux_cond_24_shl};
  assign mux_cond_25_shl = {mux_cond_25, 17'h0};
  assign mux_cond_25_pad = {2'h0,mux_cond_25_shl};
  assign mux_cond_26_shl = {mux_cond_26, 5'h0};
  assign mux_cond_26_pad = {14'h0,mux_cond_26_shl};
  assign mux_cond_27_shl = {mux_cond_27, 6'h0};
  assign mux_cond_27_pad = {13'h0,mux_cond_27_shl};
  assign mux_cond_28_shl = {mux_cond_28, 19'h0};
  assign mux_cond_28_pad = mux_cond_28_shl;
  assign mux_cond_29_shl = {mux_cond_29, 16'h0};
  assign mux_cond_29_pad = {3'h0,mux_cond_29_shl};
  assign mux_cond_30_shl = {mux_cond_30, 18'h0};
  assign mux_cond_30_pad = {1'h0,mux_cond_30_shl};
  assign mux_cond_31_shl = mux_cond_31;
  assign mux_cond_31_pad = {19'h0,mux_cond_31_shl};
  assign mux_cond_32_shl = {mux_cond_32, 2'h0};
  assign mux_cond_32_pad = {17'h0,mux_cond_32_shl};
  assign mux_cond_33_shl = {mux_cond_33, 11'h0};
  assign mux_cond_33_pad = {8'h0,mux_cond_33_shl};
  assign mux_cond_34_shl = {mux_cond_34, 18'h0};
  assign mux_cond_34_pad = {1'h0,mux_cond_34_shl};
  assign mux_cond_35_shl = {mux_cond_35, 9'h0};
  assign mux_cond_35_pad = {10'h0,mux_cond_35_shl};
  assign mux_cond_36_shl = {mux_cond_36, 1'h0};
  assign mux_cond_36_pad = {18'h0,mux_cond_36_shl};
  assign mux_cond_37_shl = {mux_cond_37, 1'h0};
  assign mux_cond_37_pad = {18'h0,mux_cond_37_shl};
  assign mux_cond_38_shl = {mux_cond_38, 3'h0};
  assign mux_cond_38_pad = {16'h0,mux_cond_38_shl};
  assign mux_cond_39_shl = mux_cond_39;
  assign mux_cond_39_pad = {19'h0,mux_cond_39_shl};
  assign mux_cond_40_shl = {mux_cond_40, 15'h0};
  assign mux_cond_40_pad = {4'h0,mux_cond_40_shl};
  assign mux_cond_41_shl = {mux_cond_41, 6'h0};
  assign mux_cond_41_pad = {13'h0,mux_cond_41_shl};
  assign mux_cond_42_shl = {mux_cond_42, 19'h0};
  assign mux_cond_42_pad = mux_cond_42_shl;
  assign mux_cond_43_shl = {mux_cond_43, 19'h0};
  assign mux_cond_43_pad = mux_cond_43_shl;
  assign mux_cond_44_shl = {mux_cond_44, 13'h0};
  assign mux_cond_44_pad = {6'h0,mux_cond_44_shl};
  assign mux_cond_45_shl = {mux_cond_45, 1'h0};
  assign mux_cond_45_pad = {18'h0,mux_cond_45_shl};
  assign mux_cond_46_shl = {mux_cond_46, 8'h0};
  assign mux_cond_46_pad = {11'h0,mux_cond_46_shl};
  assign mux_cond_47_shl = {mux_cond_47, 17'h0};
  assign mux_cond_47_pad = {2'h0,mux_cond_47_shl};
  assign mux_cond_48_shl = {mux_cond_48, 11'h0};
  assign mux_cond_48_pad = {8'h0,mux_cond_48_shl};
  assign mux_cond_49_shl = {mux_cond_49, 3'h0};
  assign mux_cond_49_pad = {16'h0,mux_cond_49_shl};
  assign mux_cond_50_shl = {mux_cond_50, 11'h0};
  assign mux_cond_50_pad = {8'h0,mux_cond_50_shl};
  assign mux_cond_51_shl = {mux_cond_51, 14'h0};
  assign mux_cond_51_pad = {5'h0,mux_cond_51_shl};
  assign mux_cond_52_shl = {mux_cond_52, 5'h0};
  assign mux_cond_52_pad = {14'h0,mux_cond_52_shl};
  assign mux_cond_53_shl = {mux_cond_53, 3'h0};
  assign mux_cond_53_pad = {16'h0,mux_cond_53_shl};
  assign mux_cond_54_shl = {mux_cond_54, 18'h0};
  assign mux_cond_54_pad = {1'h0,mux_cond_54_shl};
  assign mux_cond_55_shl = {mux_cond_55, 9'h0};
  assign mux_cond_55_pad = {10'h0,mux_cond_55_shl};
  assign mux_cond_56_shl = {mux_cond_56, 15'h0};
  assign mux_cond_56_pad = {4'h0,mux_cond_56_shl};
  assign mux_cond_57_shl = {mux_cond_57, 17'h0};
  assign mux_cond_57_pad = {2'h0,mux_cond_57_shl};
  assign mux_cond_58_shl = {mux_cond_58, 13'h0};
  assign mux_cond_58_pad = {6'h0,mux_cond_58_shl};
  assign mux_cond_59_shl = {mux_cond_59, 12'h0};
  assign mux_cond_59_pad = {7'h0,mux_cond_59_shl};
  assign mux_cond_60_shl = {mux_cond_60, 14'h0};
  assign mux_cond_60_pad = {5'h0,mux_cond_60_shl};
  assign mux_cond_61_shl = {mux_cond_61, 9'h0};
  assign mux_cond_61_pad = {10'h0,mux_cond_61_shl};
  assign mux_cond_62_shl = {mux_cond_62, 4'h0};
  assign mux_cond_62_pad = {15'h0,mux_cond_62_shl};
  assign mux_cond_63_shl = {mux_cond_63, 6'h0};
  assign mux_cond_63_pad = {13'h0,mux_cond_63_shl};
  assign mux_cond_64_shl = {mux_cond_64, 5'h0};
  assign mux_cond_64_pad = {14'h0,mux_cond_64_shl};
  assign mux_cond_65_shl = {mux_cond_65, 9'h0};
  assign mux_cond_65_pad = {10'h0,mux_cond_65_shl};
  assign mux_cond_66_shl = mux_cond_66;
  assign mux_cond_66_pad = {19'h0,mux_cond_66_shl};
  assign mux_cond_67_shl = {mux_cond_67, 13'h0};
  assign mux_cond_67_pad = {6'h0,mux_cond_67_shl};
  assign mux_cond_68_shl = {mux_cond_68, 19'h0};
  assign mux_cond_68_pad = mux_cond_68_shl;
  assign mux_cond_69_shl = {mux_cond_69, 8'h0};
  assign mux_cond_69_pad = {11'h0,mux_cond_69_shl};
  assign mux_cond_70_shl = {mux_cond_70, 7'h0};
  assign mux_cond_70_pad = {12'h0,mux_cond_70_shl};
  assign mux_cond_71_shl = {mux_cond_71, 8'h0};
  assign mux_cond_71_pad = {11'h0,mux_cond_71_shl};
  assign mux_cond_72_shl = {mux_cond_72, 3'h0};
  assign mux_cond_72_pad = {16'h0,mux_cond_72_shl};
  assign mux_cond_73_shl = {mux_cond_73, 6'h0};
  assign mux_cond_73_pad = {13'h0,mux_cond_73_shl};
  assign mux_cond_74_shl = {mux_cond_74, 18'h0};
  assign mux_cond_74_pad = {1'h0,mux_cond_74_shl};
  assign mux_cond_75_shl = {mux_cond_75, 18'h0};
  assign mux_cond_75_pad = {1'h0,mux_cond_75_shl};
  assign mux_cond_76_shl = {mux_cond_76, 6'h0};
  assign mux_cond_76_pad = {13'h0,mux_cond_76_shl};
  assign mux_cond_77_shl = {mux_cond_77, 5'h0};
  assign mux_cond_77_pad = {14'h0,mux_cond_77_shl};
  assign mux_cond_78_shl = {mux_cond_78, 14'h0};
  assign mux_cond_78_pad = {5'h0,mux_cond_78_shl};
  assign mux_cond_79_shl = {mux_cond_79, 9'h0};
  assign mux_cond_79_pad = {10'h0,mux_cond_79_shl};
  assign mux_cond_80_shl = {mux_cond_80, 8'h0};
  assign mux_cond_80_pad = {11'h0,mux_cond_80_shl};
  assign mux_cond_81_shl = {mux_cond_81, 10'h0};
  assign mux_cond_81_pad = {9'h0,mux_cond_81_shl};
  assign mux_cond_82_shl = {mux_cond_82, 2'h0};
  assign mux_cond_82_pad = {17'h0,mux_cond_82_shl};
  assign mux_cond_83_shl = {mux_cond_83, 15'h0};
  assign mux_cond_83_pad = {4'h0,mux_cond_83_shl};
  assign mux_cond_84_shl = mux_cond_84;
  assign mux_cond_84_pad = {19'h0,mux_cond_84_shl};
  assign mux_cond_85_shl = {mux_cond_85, 1'h0};
  assign mux_cond_85_pad = {18'h0,mux_cond_85_shl};
  assign mux_cond_86_shl = {mux_cond_86, 17'h0};
  assign mux_cond_86_pad = {2'h0,mux_cond_86_shl};
  assign mux_cond_87_shl = {mux_cond_87, 15'h0};
  assign mux_cond_87_pad = {4'h0,mux_cond_87_shl};
  assign mux_cond_88_shl = {mux_cond_88, 14'h0};
  assign mux_cond_88_pad = {5'h0,mux_cond_88_shl};
  assign mux_cond_89_shl = {mux_cond_89, 15'h0};
  assign mux_cond_89_pad = {4'h0,mux_cond_89_shl};
  assign mux_cond_90_shl = mux_cond_90;
  assign mux_cond_90_pad = {19'h0,mux_cond_90_shl};
  assign mux_cond_91_shl = {mux_cond_91, 5'h0};
  assign mux_cond_91_pad = {14'h0,mux_cond_91_shl};
  assign mux_cond_92_shl = {mux_cond_92, 19'h0};
  assign mux_cond_92_pad = mux_cond_92_shl;
  assign mux_cond_93_shl = {mux_cond_93, 1'h0};
  assign mux_cond_93_pad = {18'h0,mux_cond_93_shl};
  assign mux_cond_94_shl = {mux_cond_94, 11'h0};
  assign mux_cond_94_pad = {8'h0,mux_cond_94_shl};
  assign mux_cond_95_shl = {mux_cond_95, 8'h0};
  assign mux_cond_95_pad = {11'h0,mux_cond_95_shl};
  assign mux_cond_96_shl = {mux_cond_96, 16'h0};
  assign mux_cond_96_pad = {3'h0,mux_cond_96_shl};
  assign mux_cond_97_shl = {mux_cond_97, 14'h0};
  assign mux_cond_97_pad = {5'h0,mux_cond_97_shl};
  assign MulDiv_xor64 = state_pad ^ req_dw_pad;
  assign MulDiv_xor31 = resHi_pad ^ MulDiv_xor64;
  assign MulDiv_xor66 = isHi_pad ^ mux_cond_0_pad;
  assign MulDiv_xor32 = neg_out_pad ^ MulDiv_xor66;
  assign MulDiv_xor15 = MulDiv_xor31 ^ MulDiv_xor32;
  assign MulDiv_xor68 = mux_cond_2_pad ^ mux_cond_3_pad;
  assign MulDiv_xor33 = mux_cond_1_pad ^ MulDiv_xor68;
  assign MulDiv_xor70 = mux_cond_5_pad ^ mux_cond_6_pad;
  assign MulDiv_xor34 = mux_cond_4_pad ^ MulDiv_xor70;
  assign MulDiv_xor16 = MulDiv_xor33 ^ MulDiv_xor34;
  assign MulDiv_xor7 = MulDiv_xor15 ^ MulDiv_xor16;
  assign MulDiv_xor72 = mux_cond_8_pad ^ mux_cond_9_pad;
  assign MulDiv_xor35 = mux_cond_7_pad ^ MulDiv_xor72;
  assign MulDiv_xor74 = mux_cond_11_pad ^ mux_cond_12_pad;
  assign MulDiv_xor36 = mux_cond_10_pad ^ MulDiv_xor74;
  assign MulDiv_xor17 = MulDiv_xor35 ^ MulDiv_xor36;
  assign MulDiv_xor76 = mux_cond_14_pad ^ mux_cond_15_pad;
  assign MulDiv_xor37 = mux_cond_13_pad ^ MulDiv_xor76;
  assign MulDiv_xor77 = mux_cond_16_pad ^ mux_cond_17_pad;
  assign MulDiv_xor78 = mux_cond_18_pad ^ mux_cond_19_pad;
  assign MulDiv_xor38 = MulDiv_xor77 ^ MulDiv_xor78;
  assign MulDiv_xor18 = MulDiv_xor37 ^ MulDiv_xor38;
  assign MulDiv_xor8 = MulDiv_xor17 ^ MulDiv_xor18;
  assign MulDiv_xor3 = MulDiv_xor7 ^ MulDiv_xor8;
  assign MulDiv_xor80 = mux_cond_21_pad ^ mux_cond_22_pad;
  assign MulDiv_xor39 = mux_cond_20_pad ^ MulDiv_xor80;
  assign MulDiv_xor82 = mux_cond_24_pad ^ mux_cond_25_pad;
  assign MulDiv_xor40 = mux_cond_23_pad ^ MulDiv_xor82;
  assign MulDiv_xor19 = MulDiv_xor39 ^ MulDiv_xor40;
  assign MulDiv_xor84 = mux_cond_27_pad ^ mux_cond_28_pad;
  assign MulDiv_xor41 = mux_cond_26_pad ^ MulDiv_xor84;
  assign MulDiv_xor85 = mux_cond_29_pad ^ mux_cond_30_pad;
  assign MulDiv_xor86 = mux_cond_31_pad ^ mux_cond_32_pad;
  assign MulDiv_xor42 = MulDiv_xor85 ^ MulDiv_xor86;
  assign MulDiv_xor20 = MulDiv_xor41 ^ MulDiv_xor42;
  assign MulDiv_xor9 = MulDiv_xor19 ^ MulDiv_xor20;
  assign MulDiv_xor88 = mux_cond_34_pad ^ mux_cond_35_pad;
  assign MulDiv_xor43 = mux_cond_33_pad ^ MulDiv_xor88;
  assign MulDiv_xor90 = mux_cond_37_pad ^ mux_cond_38_pad;
  assign MulDiv_xor44 = mux_cond_36_pad ^ MulDiv_xor90;
  assign MulDiv_xor21 = MulDiv_xor43 ^ MulDiv_xor44;
  assign MulDiv_xor92 = mux_cond_40_pad ^ mux_cond_41_pad;
  assign MulDiv_xor45 = mux_cond_39_pad ^ MulDiv_xor92;
  assign MulDiv_xor93 = mux_cond_42_pad ^ mux_cond_43_pad;
  assign MulDiv_xor94 = mux_cond_44_pad ^ mux_cond_45_pad;
  assign MulDiv_xor46 = MulDiv_xor93 ^ MulDiv_xor94;
  assign MulDiv_xor22 = MulDiv_xor45 ^ MulDiv_xor46;
  assign MulDiv_xor10 = MulDiv_xor21 ^ MulDiv_xor22;
  assign MulDiv_xor4 = MulDiv_xor9 ^ MulDiv_xor10;
  assign MulDiv_xor1 = MulDiv_xor3 ^ MulDiv_xor4;
  assign MulDiv_xor96 = mux_cond_47_pad ^ mux_cond_48_pad;
  assign MulDiv_xor47 = mux_cond_46_pad ^ MulDiv_xor96;
  assign MulDiv_xor98 = mux_cond_50_pad ^ mux_cond_51_pad;
  assign MulDiv_xor48 = mux_cond_49_pad ^ MulDiv_xor98;
  assign MulDiv_xor23 = MulDiv_xor47 ^ MulDiv_xor48;
  assign MulDiv_xor100 = mux_cond_53_pad ^ mux_cond_54_pad;
  assign MulDiv_xor49 = mux_cond_52_pad ^ MulDiv_xor100;
  assign MulDiv_xor101 = mux_cond_55_pad ^ mux_cond_56_pad;
  assign MulDiv_xor102 = mux_cond_57_pad ^ mux_cond_58_pad;
  assign MulDiv_xor50 = MulDiv_xor101 ^ MulDiv_xor102;
  assign MulDiv_xor24 = MulDiv_xor49 ^ MulDiv_xor50;
  assign MulDiv_xor11 = MulDiv_xor23 ^ MulDiv_xor24;
  assign MulDiv_xor104 = mux_cond_60_pad ^ mux_cond_61_pad;
  assign MulDiv_xor51 = mux_cond_59_pad ^ MulDiv_xor104;
  assign MulDiv_xor106 = mux_cond_63_pad ^ mux_cond_64_pad;
  assign MulDiv_xor52 = mux_cond_62_pad ^ MulDiv_xor106;
  assign MulDiv_xor25 = MulDiv_xor51 ^ MulDiv_xor52;
  assign MulDiv_xor108 = mux_cond_66_pad ^ mux_cond_67_pad;
  assign MulDiv_xor53 = mux_cond_65_pad ^ MulDiv_xor108;
  assign MulDiv_xor109 = mux_cond_68_pad ^ mux_cond_69_pad;
  assign MulDiv_xor110 = mux_cond_70_pad ^ mux_cond_71_pad;
  assign MulDiv_xor54 = MulDiv_xor109 ^ MulDiv_xor110;
  assign MulDiv_xor26 = MulDiv_xor53 ^ MulDiv_xor54;
  assign MulDiv_xor12 = MulDiv_xor25 ^ MulDiv_xor26;
  assign MulDiv_xor5 = MulDiv_xor11 ^ MulDiv_xor12;
  assign MulDiv_xor112 = mux_cond_73_pad ^ mux_cond_74_pad;
  assign MulDiv_xor55 = mux_cond_72_pad ^ MulDiv_xor112;
  assign MulDiv_xor114 = mux_cond_76_pad ^ mux_cond_77_pad;
  assign MulDiv_xor56 = mux_cond_75_pad ^ MulDiv_xor114;
  assign MulDiv_xor27 = MulDiv_xor55 ^ MulDiv_xor56;
  assign MulDiv_xor116 = mux_cond_79_pad ^ mux_cond_80_pad;
  assign MulDiv_xor57 = mux_cond_78_pad ^ MulDiv_xor116;
  assign MulDiv_xor117 = mux_cond_81_pad ^ mux_cond_82_pad;
  assign MulDiv_xor118 = mux_cond_83_pad ^ mux_cond_84_pad;
  assign MulDiv_xor58 = MulDiv_xor117 ^ MulDiv_xor118;
  assign MulDiv_xor28 = MulDiv_xor57 ^ MulDiv_xor58;
  assign MulDiv_xor13 = MulDiv_xor27 ^ MulDiv_xor28;
  assign MulDiv_xor120 = mux_cond_86_pad ^ mux_cond_87_pad;
  assign MulDiv_xor59 = mux_cond_85_pad ^ MulDiv_xor120;
  assign MulDiv_xor122 = mux_cond_89_pad ^ mux_cond_90_pad;
  assign MulDiv_xor60 = mux_cond_88_pad ^ MulDiv_xor122;
  assign MulDiv_xor29 = MulDiv_xor59 ^ MulDiv_xor60;
  assign MulDiv_xor124 = mux_cond_92_pad ^ mux_cond_93_pad;
  assign MulDiv_xor61 = mux_cond_91_pad ^ MulDiv_xor124;
  assign MulDiv_xor125 = mux_cond_94_pad ^ mux_cond_95_pad;
  assign MulDiv_xor126 = mux_cond_96_pad ^ mux_cond_97_pad;
  assign MulDiv_xor62 = MulDiv_xor125 ^ MulDiv_xor126;
  assign MulDiv_xor30 = MulDiv_xor61 ^ MulDiv_xor62;
  assign MulDiv_xor14 = MulDiv_xor29 ^ MulDiv_xor30;
  assign MulDiv_xor6 = MulDiv_xor13 ^ MulDiv_xor14;
  assign MulDiv_xor2 = MulDiv_xor5 ^ MulDiv_xor6;
  assign MulDiv_xor0 = MulDiv_xor1 ^ MulDiv_xor2;
  assign io_covSum = MulDiv_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  req_dw = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  req_tag = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  count = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  neg_out = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  isHi = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  resHi = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {3{`RANDOM}};
  divisor = _RAND_7[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {5{`RANDOM}};
  remainder = _RAND_8[129:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  MulDiv_state = _RAND_9[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    MulDiv_cov[initvar] = _RAND_10[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  MulDiv_covSum = _RAND_11[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      state <= 3'h0;
    end else if (reset) begin
      state <= 3'h0;
    end else if (_T_474) begin
      if (cmdMul) begin
        state <= 3'h2;
      end else if (_T_475) begin
        state <= 3'h1;
      end else begin
        state <= 3'h3;
      end
    end else if (_T_473) begin
      state <= 3'h0;
    end else if (_T_125) begin
      if (_T_134) begin
        if (neg_out) begin
          state <= 3'h5;
        end else begin
          state <= 3'h7;
        end
      end else if (_T_72) begin
        if (_T_124) begin
          state <= 3'h6;
        end else if (_T_71) begin
          state <= 3'h7;
        end else if (_T_68) begin
          state <= 3'h3;
        end
      end else if (_T_71) begin
        state <= 3'h7;
      end else if (_T_68) begin
        state <= 3'h3;
      end
    end else if (_T_72) begin
      if (_T_124) begin
        state <= 3'h6;
      end else if (_T_71) begin
        state <= 3'h7;
      end else if (_T_68) begin
        state <= 3'h3;
      end
    end else if (_T_71) begin
      state <= 3'h7;
    end else if (_T_68) begin
      state <= 3'h3;
    end
    if (metaReset) begin
      req_dw <= 1'h0;
    end else if (_T_474) begin
      req_dw <= io_req_bits_dw;
    end
    if (metaReset) begin
      req_tag <= 5'h0;
    end else if (_T_474) begin
      req_tag <= io_req_bits_tag;
    end
    if (metaReset) begin
      count <= 7'h0;
    end else if (_T_474) begin
      count <= {{4'd0}, _T_481};
    end else if (_T_125) begin
      if (_T_466) begin
        count <= {{1'd0}, ~_T_460};
      end else begin
        count <= _T_122;
      end
    end else if (_T_72) begin
      count <= _T_122;
    end
    if (metaReset) begin
      neg_out <= 1'h0;
    end else if (_T_474) begin
      if (cmdHi) begin
        neg_out <= lhs_sign;
      end else begin
        neg_out <= _T_482;
      end
    end else if (_T_125) begin
      if (_T_471) begin
        neg_out <= 1'h0;
      end
    end
    if (metaReset) begin
      isHi <= 1'h0;
    end else if (_T_474) begin
      isHi <= cmdHi;
    end
    if (metaReset) begin
      resHi <= 1'h0;
    end else if (_T_474) begin
      resHi <= 1'h0;
    end else if (_T_125) begin
      if (_T_134) begin
        resHi <= isHi;
      end else if (_T_72) begin
        if (_T_124) begin
          resHi <= isHi;
        end else if (_T_71) begin
          resHi <= 1'h0;
        end
      end else if (_T_71) begin
        resHi <= 1'h0;
      end
    end else if (_T_72) begin
      if (_T_124) begin
        resHi <= isHi;
      end else if (_T_71) begin
        resHi <= 1'h0;
      end
    end else if (_T_71) begin
      resHi <= 1'h0;
    end
    if (metaReset) begin
      divisor <= 65'h0;
    end else if (_T_474) begin
      divisor <= _T_484;
    end else if (_T_68) begin
      if (divisor[63]) begin
        divisor <= subtractor;
      end
    end
    if (metaReset) begin
      remainder <= 130'h0;
    end else if (_T_474) begin
      remainder <= {{66'd0}, lhs_in};
    end else if (_T_125) begin
      remainder <= {{1'd0}, _GEN_16};
    end else if (_T_72) begin
      remainder <= _T_120;
    end else if (_T_71) begin
      remainder <= {{66'd0}, negated_remainder};
    end else if (_T_68) begin
      if (remainder[63]) begin
        remainder <= {{66'd0}, negated_remainder};
      end
    end
    MulDiv_state <= MulDiv_xor0;
    if (!(MulDiv_cov_read_data)) begin
      MulDiv_covSum <= MulDiv_covSum + 1'h1;
    end
  end
  always @(posedge clock) begin
    if(MulDiv_cov_write_en & MulDiv_cov_write_mask) begin
      MulDiv_cov[MulDiv_cov_write_addr] <= MulDiv_cov_write_data; // @[Coverage map for MulDiv]
    end
  end
endmodule
module PMPChecker(
  input  [1:0]  io_prv,
  input         io_pmp_0_cfg_l,
  input  [1:0]  io_pmp_0_cfg_a,
  input         io_pmp_0_cfg_x,
  input         io_pmp_0_cfg_w,
  input         io_pmp_0_cfg_r,
  input  [29:0] io_pmp_0_addr,
  input  [31:0] io_pmp_0_mask,
  input         io_pmp_1_cfg_l,
  input  [1:0]  io_pmp_1_cfg_a,
  input         io_pmp_1_cfg_x,
  input         io_pmp_1_cfg_w,
  input         io_pmp_1_cfg_r,
  input  [29:0] io_pmp_1_addr,
  input  [31:0] io_pmp_1_mask,
  input         io_pmp_2_cfg_l,
  input  [1:0]  io_pmp_2_cfg_a,
  input         io_pmp_2_cfg_x,
  input         io_pmp_2_cfg_w,
  input         io_pmp_2_cfg_r,
  input  [29:0] io_pmp_2_addr,
  input  [31:0] io_pmp_2_mask,
  input         io_pmp_3_cfg_l,
  input  [1:0]  io_pmp_3_cfg_a,
  input         io_pmp_3_cfg_x,
  input         io_pmp_3_cfg_w,
  input         io_pmp_3_cfg_r,
  input  [29:0] io_pmp_3_addr,
  input  [31:0] io_pmp_3_mask,
  input         io_pmp_4_cfg_l,
  input  [1:0]  io_pmp_4_cfg_a,
  input         io_pmp_4_cfg_x,
  input         io_pmp_4_cfg_w,
  input         io_pmp_4_cfg_r,
  input  [29:0] io_pmp_4_addr,
  input  [31:0] io_pmp_4_mask,
  input         io_pmp_5_cfg_l,
  input  [1:0]  io_pmp_5_cfg_a,
  input         io_pmp_5_cfg_x,
  input         io_pmp_5_cfg_w,
  input         io_pmp_5_cfg_r,
  input  [29:0] io_pmp_5_addr,
  input  [31:0] io_pmp_5_mask,
  input         io_pmp_6_cfg_l,
  input  [1:0]  io_pmp_6_cfg_a,
  input         io_pmp_6_cfg_x,
  input         io_pmp_6_cfg_w,
  input         io_pmp_6_cfg_r,
  input  [29:0] io_pmp_6_addr,
  input  [31:0] io_pmp_6_mask,
  input         io_pmp_7_cfg_l,
  input  [1:0]  io_pmp_7_cfg_a,
  input         io_pmp_7_cfg_x,
  input         io_pmp_7_cfg_w,
  input         io_pmp_7_cfg_r,
  input  [29:0] io_pmp_7_addr,
  input  [31:0] io_pmp_7_mask,
  input  [31:0] io_addr,
  input  [1:0]  io_size,
  output        io_r,
  output        io_w,
  output        io_x,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  default_; // @[PMP.scala 149:56]
  wire [5:0] _T_39; // @[package.scala 185:77]
  wire [31:0] _GEN_0; // @[PMP.scala 62:26]
  wire [31:0] _T_42; // @[PMP.scala 62:26]
  wire [31:0] _T_44; // @[PMP.scala 54:36]
  wire [31:0] _T_46; // @[PMP.scala 54:48]
  wire [28:0] _T_48; // @[PMP.scala 63:53]
  wire [28:0] _T_50; // @[PMP.scala 57:47]
  wire [28:0] _T_52; // @[PMP.scala 57:52]
  wire  _T_53; // @[PMP.scala 57:58]
  wire [2:0] _T_59; // @[PMP.scala 64:55]
  wire [2:0] _T_61; // @[PMP.scala 57:47]
  wire [2:0] _T_63; // @[PMP.scala 57:52]
  wire  _T_64; // @[PMP.scala 57:58]
  wire  _T_65; // @[PMP.scala 65:16]
  wire [31:0] _T_72; // @[PMP.scala 54:36]
  wire [31:0] _T_74; // @[PMP.scala 54:48]
  wire [28:0] _T_76; // @[PMP.scala 74:52]
  wire  _T_77; // @[PMP.scala 74:39]
  wire [28:0] _T_84; // @[PMP.scala 75:41]
  wire  _T_85; // @[PMP.scala 75:69]
  wire [2:0] _T_87; // @[PMP.scala 76:42]
  wire [2:0] _T_92; // @[PMP.scala 76:64]
  wire  _T_93; // @[PMP.scala 76:53]
  wire  _T_94; // @[PMP.scala 77:30]
  wire  _T_95; // @[PMP.scala 77:16]
  wire  _T_103; // @[PMP.scala 74:39]
  wire  _T_111; // @[PMP.scala 75:69]
  wire  _T_119; // @[PMP.scala 76:53]
  wire  _T_120; // @[PMP.scala 77:30]
  wire  _T_121; // @[PMP.scala 77:16]
  wire  _T_122; // @[PMP.scala 88:48]
  wire  _T_123; // @[PMP.scala 126:61]
  wire  _T_124; // @[PMP.scala 126:8]
  wire  _T_126; // @[PMP.scala 157:26]
  wire [2:0] _T_146; // @[PMP.scala 117:123]
  wire  _T_147; // @[PMP.scala 117:145]
  wire  _T_148; // @[PMP.scala 117:88]
  wire [2:0] _T_164; // @[PMP.scala 118:113]
  wire  _T_165; // @[PMP.scala 118:146]
  wire  _T_166; // @[PMP.scala 118:83]
  wire  _T_167; // @[PMP.scala 119:46]
  wire [2:0] _T_171; // @[PMP.scala 120:32]
  wire  _T_172; // @[PMP.scala 120:57]
  wire  _T_174; // @[PMP.scala 121:8]
  wire  _T_177; // @[PMP.scala 160:27]
  wire  _T_178; // @[PMP.scala 160:41]
  wire  _T_179; // @[PMP.scala 161:27]
  wire  _T_180; // @[PMP.scala 161:41]
  wire  _T_181; // @[PMP.scala 162:27]
  wire  _T_182; // @[PMP.scala 162:41]
  wire  _T_183_cfg_x; // @[PMP.scala 163:8]
  wire  _T_183_cfg_w; // @[PMP.scala 163:8]
  wire  _T_183_cfg_r; // @[PMP.scala 163:8]
  wire [31:0] _T_189; // @[PMP.scala 62:26]
  wire [28:0] _T_199; // @[PMP.scala 57:52]
  wire  _T_200; // @[PMP.scala 57:58]
  wire [2:0] _T_208; // @[PMP.scala 57:47]
  wire [2:0] _T_210; // @[PMP.scala 57:52]
  wire  _T_211; // @[PMP.scala 57:58]
  wire  _T_212; // @[PMP.scala 65:16]
  wire [31:0] _T_219; // @[PMP.scala 54:36]
  wire [31:0] _T_221; // @[PMP.scala 54:48]
  wire [28:0] _T_223; // @[PMP.scala 74:52]
  wire  _T_224; // @[PMP.scala 74:39]
  wire [28:0] _T_231; // @[PMP.scala 75:41]
  wire  _T_232; // @[PMP.scala 75:69]
  wire [2:0] _T_239; // @[PMP.scala 76:64]
  wire  _T_240; // @[PMP.scala 76:53]
  wire  _T_241; // @[PMP.scala 77:30]
  wire  _T_242; // @[PMP.scala 77:16]
  wire  _T_266; // @[PMP.scala 76:53]
  wire  _T_267; // @[PMP.scala 77:30]
  wire  _T_268; // @[PMP.scala 77:16]
  wire  _T_269; // @[PMP.scala 88:48]
  wire  _T_270; // @[PMP.scala 126:61]
  wire  _T_271; // @[PMP.scala 126:8]
  wire  _T_273; // @[PMP.scala 157:26]
  wire [2:0] _T_293; // @[PMP.scala 117:123]
  wire  _T_294; // @[PMP.scala 117:145]
  wire  _T_295; // @[PMP.scala 117:88]
  wire [2:0] _T_311; // @[PMP.scala 118:113]
  wire  _T_312; // @[PMP.scala 118:146]
  wire  _T_313; // @[PMP.scala 118:83]
  wire  _T_314; // @[PMP.scala 119:46]
  wire [2:0] _T_318; // @[PMP.scala 120:32]
  wire  _T_319; // @[PMP.scala 120:57]
  wire  _T_321; // @[PMP.scala 121:8]
  wire  _T_324; // @[PMP.scala 160:27]
  wire  _T_325; // @[PMP.scala 160:41]
  wire  _T_326; // @[PMP.scala 161:27]
  wire  _T_327; // @[PMP.scala 161:41]
  wire  _T_328; // @[PMP.scala 162:27]
  wire  _T_329; // @[PMP.scala 162:41]
  wire  _T_330_cfg_x; // @[PMP.scala 163:8]
  wire  _T_330_cfg_w; // @[PMP.scala 163:8]
  wire  _T_330_cfg_r; // @[PMP.scala 163:8]
  wire [31:0] _T_336; // @[PMP.scala 62:26]
  wire [28:0] _T_346; // @[PMP.scala 57:52]
  wire  _T_347; // @[PMP.scala 57:58]
  wire [2:0] _T_355; // @[PMP.scala 57:47]
  wire [2:0] _T_357; // @[PMP.scala 57:52]
  wire  _T_358; // @[PMP.scala 57:58]
  wire  _T_359; // @[PMP.scala 65:16]
  wire [31:0] _T_366; // @[PMP.scala 54:36]
  wire [31:0] _T_368; // @[PMP.scala 54:48]
  wire [28:0] _T_370; // @[PMP.scala 74:52]
  wire  _T_371; // @[PMP.scala 74:39]
  wire [28:0] _T_378; // @[PMP.scala 75:41]
  wire  _T_379; // @[PMP.scala 75:69]
  wire [2:0] _T_386; // @[PMP.scala 76:64]
  wire  _T_387; // @[PMP.scala 76:53]
  wire  _T_388; // @[PMP.scala 77:30]
  wire  _T_389; // @[PMP.scala 77:16]
  wire  _T_413; // @[PMP.scala 76:53]
  wire  _T_414; // @[PMP.scala 77:30]
  wire  _T_415; // @[PMP.scala 77:16]
  wire  _T_416; // @[PMP.scala 88:48]
  wire  _T_417; // @[PMP.scala 126:61]
  wire  _T_418; // @[PMP.scala 126:8]
  wire  _T_420; // @[PMP.scala 157:26]
  wire [2:0] _T_440; // @[PMP.scala 117:123]
  wire  _T_441; // @[PMP.scala 117:145]
  wire  _T_442; // @[PMP.scala 117:88]
  wire [2:0] _T_458; // @[PMP.scala 118:113]
  wire  _T_459; // @[PMP.scala 118:146]
  wire  _T_460; // @[PMP.scala 118:83]
  wire  _T_461; // @[PMP.scala 119:46]
  wire [2:0] _T_465; // @[PMP.scala 120:32]
  wire  _T_466; // @[PMP.scala 120:57]
  wire  _T_468; // @[PMP.scala 121:8]
  wire  _T_471; // @[PMP.scala 160:27]
  wire  _T_472; // @[PMP.scala 160:41]
  wire  _T_473; // @[PMP.scala 161:27]
  wire  _T_474; // @[PMP.scala 161:41]
  wire  _T_475; // @[PMP.scala 162:27]
  wire  _T_476; // @[PMP.scala 162:41]
  wire  _T_477_cfg_x; // @[PMP.scala 163:8]
  wire  _T_477_cfg_w; // @[PMP.scala 163:8]
  wire  _T_477_cfg_r; // @[PMP.scala 163:8]
  wire [31:0] _T_483; // @[PMP.scala 62:26]
  wire [28:0] _T_493; // @[PMP.scala 57:52]
  wire  _T_494; // @[PMP.scala 57:58]
  wire [2:0] _T_502; // @[PMP.scala 57:47]
  wire [2:0] _T_504; // @[PMP.scala 57:52]
  wire  _T_505; // @[PMP.scala 57:58]
  wire  _T_506; // @[PMP.scala 65:16]
  wire [31:0] _T_513; // @[PMP.scala 54:36]
  wire [31:0] _T_515; // @[PMP.scala 54:48]
  wire [28:0] _T_517; // @[PMP.scala 74:52]
  wire  _T_518; // @[PMP.scala 74:39]
  wire [28:0] _T_525; // @[PMP.scala 75:41]
  wire  _T_526; // @[PMP.scala 75:69]
  wire [2:0] _T_533; // @[PMP.scala 76:64]
  wire  _T_534; // @[PMP.scala 76:53]
  wire  _T_535; // @[PMP.scala 77:30]
  wire  _T_536; // @[PMP.scala 77:16]
  wire  _T_560; // @[PMP.scala 76:53]
  wire  _T_561; // @[PMP.scala 77:30]
  wire  _T_562; // @[PMP.scala 77:16]
  wire  _T_563; // @[PMP.scala 88:48]
  wire  _T_564; // @[PMP.scala 126:61]
  wire  _T_565; // @[PMP.scala 126:8]
  wire  _T_567; // @[PMP.scala 157:26]
  wire [2:0] _T_587; // @[PMP.scala 117:123]
  wire  _T_588; // @[PMP.scala 117:145]
  wire  _T_589; // @[PMP.scala 117:88]
  wire [2:0] _T_605; // @[PMP.scala 118:113]
  wire  _T_606; // @[PMP.scala 118:146]
  wire  _T_607; // @[PMP.scala 118:83]
  wire  _T_608; // @[PMP.scala 119:46]
  wire [2:0] _T_612; // @[PMP.scala 120:32]
  wire  _T_613; // @[PMP.scala 120:57]
  wire  _T_615; // @[PMP.scala 121:8]
  wire  _T_618; // @[PMP.scala 160:27]
  wire  _T_619; // @[PMP.scala 160:41]
  wire  _T_620; // @[PMP.scala 161:27]
  wire  _T_621; // @[PMP.scala 161:41]
  wire  _T_622; // @[PMP.scala 162:27]
  wire  _T_623; // @[PMP.scala 162:41]
  wire  _T_624_cfg_x; // @[PMP.scala 163:8]
  wire  _T_624_cfg_w; // @[PMP.scala 163:8]
  wire  _T_624_cfg_r; // @[PMP.scala 163:8]
  wire [31:0] _T_630; // @[PMP.scala 62:26]
  wire [28:0] _T_640; // @[PMP.scala 57:52]
  wire  _T_641; // @[PMP.scala 57:58]
  wire [2:0] _T_649; // @[PMP.scala 57:47]
  wire [2:0] _T_651; // @[PMP.scala 57:52]
  wire  _T_652; // @[PMP.scala 57:58]
  wire  _T_653; // @[PMP.scala 65:16]
  wire [31:0] _T_660; // @[PMP.scala 54:36]
  wire [31:0] _T_662; // @[PMP.scala 54:48]
  wire [28:0] _T_664; // @[PMP.scala 74:52]
  wire  _T_665; // @[PMP.scala 74:39]
  wire [28:0] _T_672; // @[PMP.scala 75:41]
  wire  _T_673; // @[PMP.scala 75:69]
  wire [2:0] _T_680; // @[PMP.scala 76:64]
  wire  _T_681; // @[PMP.scala 76:53]
  wire  _T_682; // @[PMP.scala 77:30]
  wire  _T_683; // @[PMP.scala 77:16]
  wire  _T_707; // @[PMP.scala 76:53]
  wire  _T_708; // @[PMP.scala 77:30]
  wire  _T_709; // @[PMP.scala 77:16]
  wire  _T_710; // @[PMP.scala 88:48]
  wire  _T_711; // @[PMP.scala 126:61]
  wire  _T_712; // @[PMP.scala 126:8]
  wire  _T_714; // @[PMP.scala 157:26]
  wire [2:0] _T_734; // @[PMP.scala 117:123]
  wire  _T_735; // @[PMP.scala 117:145]
  wire  _T_736; // @[PMP.scala 117:88]
  wire [2:0] _T_752; // @[PMP.scala 118:113]
  wire  _T_753; // @[PMP.scala 118:146]
  wire  _T_754; // @[PMP.scala 118:83]
  wire  _T_755; // @[PMP.scala 119:46]
  wire [2:0] _T_759; // @[PMP.scala 120:32]
  wire  _T_760; // @[PMP.scala 120:57]
  wire  _T_762; // @[PMP.scala 121:8]
  wire  _T_765; // @[PMP.scala 160:27]
  wire  _T_766; // @[PMP.scala 160:41]
  wire  _T_767; // @[PMP.scala 161:27]
  wire  _T_768; // @[PMP.scala 161:41]
  wire  _T_769; // @[PMP.scala 162:27]
  wire  _T_770; // @[PMP.scala 162:41]
  wire  _T_771_cfg_x; // @[PMP.scala 163:8]
  wire  _T_771_cfg_w; // @[PMP.scala 163:8]
  wire  _T_771_cfg_r; // @[PMP.scala 163:8]
  wire [31:0] _T_777; // @[PMP.scala 62:26]
  wire [28:0] _T_787; // @[PMP.scala 57:52]
  wire  _T_788; // @[PMP.scala 57:58]
  wire [2:0] _T_796; // @[PMP.scala 57:47]
  wire [2:0] _T_798; // @[PMP.scala 57:52]
  wire  _T_799; // @[PMP.scala 57:58]
  wire  _T_800; // @[PMP.scala 65:16]
  wire [31:0] _T_807; // @[PMP.scala 54:36]
  wire [31:0] _T_809; // @[PMP.scala 54:48]
  wire [28:0] _T_811; // @[PMP.scala 74:52]
  wire  _T_812; // @[PMP.scala 74:39]
  wire [28:0] _T_819; // @[PMP.scala 75:41]
  wire  _T_820; // @[PMP.scala 75:69]
  wire [2:0] _T_827; // @[PMP.scala 76:64]
  wire  _T_828; // @[PMP.scala 76:53]
  wire  _T_829; // @[PMP.scala 77:30]
  wire  _T_830; // @[PMP.scala 77:16]
  wire  _T_854; // @[PMP.scala 76:53]
  wire  _T_855; // @[PMP.scala 77:30]
  wire  _T_856; // @[PMP.scala 77:16]
  wire  _T_857; // @[PMP.scala 88:48]
  wire  _T_858; // @[PMP.scala 126:61]
  wire  _T_859; // @[PMP.scala 126:8]
  wire  _T_861; // @[PMP.scala 157:26]
  wire [2:0] _T_881; // @[PMP.scala 117:123]
  wire  _T_882; // @[PMP.scala 117:145]
  wire  _T_883; // @[PMP.scala 117:88]
  wire [2:0] _T_899; // @[PMP.scala 118:113]
  wire  _T_900; // @[PMP.scala 118:146]
  wire  _T_901; // @[PMP.scala 118:83]
  wire  _T_902; // @[PMP.scala 119:46]
  wire [2:0] _T_906; // @[PMP.scala 120:32]
  wire  _T_907; // @[PMP.scala 120:57]
  wire  _T_909; // @[PMP.scala 121:8]
  wire  _T_912; // @[PMP.scala 160:27]
  wire  _T_913; // @[PMP.scala 160:41]
  wire  _T_914; // @[PMP.scala 161:27]
  wire  _T_915; // @[PMP.scala 161:41]
  wire  _T_916; // @[PMP.scala 162:27]
  wire  _T_917; // @[PMP.scala 162:41]
  wire  _T_918_cfg_x; // @[PMP.scala 163:8]
  wire  _T_918_cfg_w; // @[PMP.scala 163:8]
  wire  _T_918_cfg_r; // @[PMP.scala 163:8]
  wire [31:0] _T_924; // @[PMP.scala 62:26]
  wire [28:0] _T_934; // @[PMP.scala 57:52]
  wire  _T_935; // @[PMP.scala 57:58]
  wire [2:0] _T_943; // @[PMP.scala 57:47]
  wire [2:0] _T_945; // @[PMP.scala 57:52]
  wire  _T_946; // @[PMP.scala 57:58]
  wire  _T_947; // @[PMP.scala 65:16]
  wire [31:0] _T_954; // @[PMP.scala 54:36]
  wire [31:0] _T_956; // @[PMP.scala 54:48]
  wire [28:0] _T_958; // @[PMP.scala 74:52]
  wire  _T_959; // @[PMP.scala 74:39]
  wire [28:0] _T_966; // @[PMP.scala 75:41]
  wire  _T_967; // @[PMP.scala 75:69]
  wire [2:0] _T_974; // @[PMP.scala 76:64]
  wire  _T_975; // @[PMP.scala 76:53]
  wire  _T_976; // @[PMP.scala 77:30]
  wire  _T_977; // @[PMP.scala 77:16]
  wire  _T_1001; // @[PMP.scala 76:53]
  wire  _T_1002; // @[PMP.scala 77:30]
  wire  _T_1003; // @[PMP.scala 77:16]
  wire  _T_1004; // @[PMP.scala 88:48]
  wire  _T_1005; // @[PMP.scala 126:61]
  wire  _T_1006; // @[PMP.scala 126:8]
  wire  _T_1008; // @[PMP.scala 157:26]
  wire [2:0] _T_1028; // @[PMP.scala 117:123]
  wire  _T_1029; // @[PMP.scala 117:145]
  wire  _T_1030; // @[PMP.scala 117:88]
  wire [2:0] _T_1046; // @[PMP.scala 118:113]
  wire  _T_1047; // @[PMP.scala 118:146]
  wire  _T_1048; // @[PMP.scala 118:83]
  wire  _T_1049; // @[PMP.scala 119:46]
  wire [2:0] _T_1053; // @[PMP.scala 120:32]
  wire  _T_1054; // @[PMP.scala 120:57]
  wire  _T_1056; // @[PMP.scala 121:8]
  wire  _T_1059; // @[PMP.scala 160:27]
  wire  _T_1060; // @[PMP.scala 160:41]
  wire  _T_1061; // @[PMP.scala 161:27]
  wire  _T_1062; // @[PMP.scala 161:41]
  wire  _T_1063; // @[PMP.scala 162:27]
  wire  _T_1064; // @[PMP.scala 162:41]
  wire  _T_1065_cfg_x; // @[PMP.scala 163:8]
  wire  _T_1065_cfg_w; // @[PMP.scala 163:8]
  wire  _T_1065_cfg_r; // @[PMP.scala 163:8]
  wire [31:0] _T_1071; // @[PMP.scala 62:26]
  wire [28:0] _T_1081; // @[PMP.scala 57:52]
  wire  _T_1082; // @[PMP.scala 57:58]
  wire [2:0] _T_1090; // @[PMP.scala 57:47]
  wire [2:0] _T_1092; // @[PMP.scala 57:52]
  wire  _T_1093; // @[PMP.scala 57:58]
  wire  _T_1094; // @[PMP.scala 65:16]
  wire  _T_1148; // @[PMP.scala 76:53]
  wire  _T_1149; // @[PMP.scala 77:30]
  wire  _T_1150; // @[PMP.scala 77:16]
  wire  _T_1152; // @[PMP.scala 126:61]
  wire  _T_1153; // @[PMP.scala 126:8]
  wire  _T_1155; // @[PMP.scala 157:26]
  wire [2:0] _T_1193; // @[PMP.scala 118:113]
  wire  _T_1194; // @[PMP.scala 118:146]
  wire  _T_1195; // @[PMP.scala 118:83]
  wire [2:0] _T_1200; // @[PMP.scala 120:32]
  wire  _T_1201; // @[PMP.scala 120:57]
  wire  _T_1203; // @[PMP.scala 121:8]
  wire  _T_1206; // @[PMP.scala 160:27]
  wire  _T_1207; // @[PMP.scala 160:41]
  wire  _T_1208; // @[PMP.scala 161:27]
  wire  _T_1209; // @[PMP.scala 161:41]
  wire  _T_1210; // @[PMP.scala 162:27]
  wire  _T_1211; // @[PMP.scala 162:41]
  wire [29:0] PMPChecker_covSum;
  assign default_ = io_prv > 2'h1; // @[PMP.scala 149:56]
  assign _T_39 = 6'h7 << io_size; // @[package.scala 185:77]
  assign _GEN_0 = {{29'd0}, ~_T_39[2:0]}; // @[PMP.scala 62:26]
  assign _T_42 = io_pmp_7_mask | _GEN_0; // @[PMP.scala 62:26]
  assign _T_44 = {io_pmp_7_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_46 = ~_T_44 | 32'h3; // @[PMP.scala 54:48]
  assign _T_48 = ~_T_46[31:3]; // @[PMP.scala 63:53]
  assign _T_50 = io_addr[31:3] ^ _T_48; // @[PMP.scala 57:47]
  assign _T_52 = _T_50 & ~io_pmp_7_mask[31:3]; // @[PMP.scala 57:52]
  assign _T_53 = _T_52 == 29'h0; // @[PMP.scala 57:58]
  assign _T_59 = ~_T_46[2:0]; // @[PMP.scala 64:55]
  assign _T_61 = io_addr[2:0] ^ _T_59; // @[PMP.scala 57:47]
  assign _T_63 = _T_61 & ~_T_42[2:0]; // @[PMP.scala 57:52]
  assign _T_64 = _T_63 == 3'h0; // @[PMP.scala 57:58]
  assign _T_65 = _T_53 & _T_64; // @[PMP.scala 65:16]
  assign _T_72 = {io_pmp_6_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_74 = ~_T_72 | 32'h3; // @[PMP.scala 54:48]
  assign _T_76 = ~_T_74[31:3]; // @[PMP.scala 74:52]
  assign _T_77 = io_addr[31:3] < _T_76; // @[PMP.scala 74:39]
  assign _T_84 = io_addr[31:3] ^ _T_76; // @[PMP.scala 75:41]
  assign _T_85 = _T_84 == 29'h0; // @[PMP.scala 75:69]
  assign _T_87 = io_addr[2:0] | ~_T_39[2:0]; // @[PMP.scala 76:42]
  assign _T_92 = ~_T_74[2:0]; // @[PMP.scala 76:64]
  assign _T_93 = _T_87 < _T_92; // @[PMP.scala 76:53]
  assign _T_94 = _T_85 & _T_93; // @[PMP.scala 77:30]
  assign _T_95 = _T_77 | _T_94; // @[PMP.scala 77:16]
  assign _T_103 = io_addr[31:3] < _T_48; // @[PMP.scala 74:39]
  assign _T_111 = _T_50 == 29'h0; // @[PMP.scala 75:69]
  assign _T_119 = io_addr[2:0] < _T_59; // @[PMP.scala 76:53]
  assign _T_120 = _T_111 & _T_119; // @[PMP.scala 77:30]
  assign _T_121 = _T_103 | _T_120; // @[PMP.scala 77:16]
  assign _T_122 = ~_T_95 & _T_121; // @[PMP.scala 88:48]
  assign _T_123 = io_pmp_7_cfg_a[0] & _T_122; // @[PMP.scala 126:61]
  assign _T_124 = io_pmp_7_cfg_a[1] ? _T_65 : _T_123; // @[PMP.scala 126:8]
  assign _T_126 = default_ & ~io_pmp_7_cfg_l; // @[PMP.scala 157:26]
  assign _T_146 = _T_92 & ~io_addr[2:0]; // @[PMP.scala 117:123]
  assign _T_147 = _T_146 != 3'h0; // @[PMP.scala 117:145]
  assign _T_148 = _T_85 & _T_147; // @[PMP.scala 117:88]
  assign _T_164 = _T_59 & _T_87; // @[PMP.scala 118:113]
  assign _T_165 = _T_164 != 3'h0; // @[PMP.scala 118:146]
  assign _T_166 = _T_111 & _T_165; // @[PMP.scala 118:83]
  assign _T_167 = _T_148 | _T_166; // @[PMP.scala 119:46]
  assign _T_171 = ~_T_39[2:0] & ~io_pmp_7_mask[2:0]; // @[PMP.scala 120:32]
  assign _T_172 = _T_171 == 3'h0; // @[PMP.scala 120:57]
  assign _T_174 = io_pmp_7_cfg_a[1] ? _T_172 : ~_T_167; // @[PMP.scala 121:8]
  assign _T_177 = _T_174 & io_pmp_7_cfg_r; // @[PMP.scala 160:27]
  assign _T_178 = _T_177 | _T_126; // @[PMP.scala 160:41]
  assign _T_179 = _T_174 & io_pmp_7_cfg_w; // @[PMP.scala 161:27]
  assign _T_180 = _T_179 | _T_126; // @[PMP.scala 161:41]
  assign _T_181 = _T_174 & io_pmp_7_cfg_x; // @[PMP.scala 162:27]
  assign _T_182 = _T_181 | _T_126; // @[PMP.scala 162:41]
  assign _T_183_cfg_x = _T_124 ? _T_182 : default_; // @[PMP.scala 163:8]
  assign _T_183_cfg_w = _T_124 ? _T_180 : default_; // @[PMP.scala 163:8]
  assign _T_183_cfg_r = _T_124 ? _T_178 : default_; // @[PMP.scala 163:8]
  assign _T_189 = io_pmp_6_mask | _GEN_0; // @[PMP.scala 62:26]
  assign _T_199 = _T_84 & ~io_pmp_6_mask[31:3]; // @[PMP.scala 57:52]
  assign _T_200 = _T_199 == 29'h0; // @[PMP.scala 57:58]
  assign _T_208 = io_addr[2:0] ^ _T_92; // @[PMP.scala 57:47]
  assign _T_210 = _T_208 & ~_T_189[2:0]; // @[PMP.scala 57:52]
  assign _T_211 = _T_210 == 3'h0; // @[PMP.scala 57:58]
  assign _T_212 = _T_200 & _T_211; // @[PMP.scala 65:16]
  assign _T_219 = {io_pmp_5_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_221 = ~_T_219 | 32'h3; // @[PMP.scala 54:48]
  assign _T_223 = ~_T_221[31:3]; // @[PMP.scala 74:52]
  assign _T_224 = io_addr[31:3] < _T_223; // @[PMP.scala 74:39]
  assign _T_231 = io_addr[31:3] ^ _T_223; // @[PMP.scala 75:41]
  assign _T_232 = _T_231 == 29'h0; // @[PMP.scala 75:69]
  assign _T_239 = ~_T_221[2:0]; // @[PMP.scala 76:64]
  assign _T_240 = _T_87 < _T_239; // @[PMP.scala 76:53]
  assign _T_241 = _T_232 & _T_240; // @[PMP.scala 77:30]
  assign _T_242 = _T_224 | _T_241; // @[PMP.scala 77:16]
  assign _T_266 = io_addr[2:0] < _T_92; // @[PMP.scala 76:53]
  assign _T_267 = _T_85 & _T_266; // @[PMP.scala 77:30]
  assign _T_268 = _T_77 | _T_267; // @[PMP.scala 77:16]
  assign _T_269 = ~_T_242 & _T_268; // @[PMP.scala 88:48]
  assign _T_270 = io_pmp_6_cfg_a[0] & _T_269; // @[PMP.scala 126:61]
  assign _T_271 = io_pmp_6_cfg_a[1] ? _T_212 : _T_270; // @[PMP.scala 126:8]
  assign _T_273 = default_ & ~io_pmp_6_cfg_l; // @[PMP.scala 157:26]
  assign _T_293 = _T_239 & ~io_addr[2:0]; // @[PMP.scala 117:123]
  assign _T_294 = _T_293 != 3'h0; // @[PMP.scala 117:145]
  assign _T_295 = _T_232 & _T_294; // @[PMP.scala 117:88]
  assign _T_311 = _T_92 & _T_87; // @[PMP.scala 118:113]
  assign _T_312 = _T_311 != 3'h0; // @[PMP.scala 118:146]
  assign _T_313 = _T_85 & _T_312; // @[PMP.scala 118:83]
  assign _T_314 = _T_295 | _T_313; // @[PMP.scala 119:46]
  assign _T_318 = ~_T_39[2:0] & ~io_pmp_6_mask[2:0]; // @[PMP.scala 120:32]
  assign _T_319 = _T_318 == 3'h0; // @[PMP.scala 120:57]
  assign _T_321 = io_pmp_6_cfg_a[1] ? _T_319 : ~_T_314; // @[PMP.scala 121:8]
  assign _T_324 = _T_321 & io_pmp_6_cfg_r; // @[PMP.scala 160:27]
  assign _T_325 = _T_324 | _T_273; // @[PMP.scala 160:41]
  assign _T_326 = _T_321 & io_pmp_6_cfg_w; // @[PMP.scala 161:27]
  assign _T_327 = _T_326 | _T_273; // @[PMP.scala 161:41]
  assign _T_328 = _T_321 & io_pmp_6_cfg_x; // @[PMP.scala 162:27]
  assign _T_329 = _T_328 | _T_273; // @[PMP.scala 162:41]
  assign _T_330_cfg_x = _T_271 ? _T_329 : _T_183_cfg_x; // @[PMP.scala 163:8]
  assign _T_330_cfg_w = _T_271 ? _T_327 : _T_183_cfg_w; // @[PMP.scala 163:8]
  assign _T_330_cfg_r = _T_271 ? _T_325 : _T_183_cfg_r; // @[PMP.scala 163:8]
  assign _T_336 = io_pmp_5_mask | _GEN_0; // @[PMP.scala 62:26]
  assign _T_346 = _T_231 & ~io_pmp_5_mask[31:3]; // @[PMP.scala 57:52]
  assign _T_347 = _T_346 == 29'h0; // @[PMP.scala 57:58]
  assign _T_355 = io_addr[2:0] ^ _T_239; // @[PMP.scala 57:47]
  assign _T_357 = _T_355 & ~_T_336[2:0]; // @[PMP.scala 57:52]
  assign _T_358 = _T_357 == 3'h0; // @[PMP.scala 57:58]
  assign _T_359 = _T_347 & _T_358; // @[PMP.scala 65:16]
  assign _T_366 = {io_pmp_4_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_368 = ~_T_366 | 32'h3; // @[PMP.scala 54:48]
  assign _T_370 = ~_T_368[31:3]; // @[PMP.scala 74:52]
  assign _T_371 = io_addr[31:3] < _T_370; // @[PMP.scala 74:39]
  assign _T_378 = io_addr[31:3] ^ _T_370; // @[PMP.scala 75:41]
  assign _T_379 = _T_378 == 29'h0; // @[PMP.scala 75:69]
  assign _T_386 = ~_T_368[2:0]; // @[PMP.scala 76:64]
  assign _T_387 = _T_87 < _T_386; // @[PMP.scala 76:53]
  assign _T_388 = _T_379 & _T_387; // @[PMP.scala 77:30]
  assign _T_389 = _T_371 | _T_388; // @[PMP.scala 77:16]
  assign _T_413 = io_addr[2:0] < _T_239; // @[PMP.scala 76:53]
  assign _T_414 = _T_232 & _T_413; // @[PMP.scala 77:30]
  assign _T_415 = _T_224 | _T_414; // @[PMP.scala 77:16]
  assign _T_416 = ~_T_389 & _T_415; // @[PMP.scala 88:48]
  assign _T_417 = io_pmp_5_cfg_a[0] & _T_416; // @[PMP.scala 126:61]
  assign _T_418 = io_pmp_5_cfg_a[1] ? _T_359 : _T_417; // @[PMP.scala 126:8]
  assign _T_420 = default_ & ~io_pmp_5_cfg_l; // @[PMP.scala 157:26]
  assign _T_440 = _T_386 & ~io_addr[2:0]; // @[PMP.scala 117:123]
  assign _T_441 = _T_440 != 3'h0; // @[PMP.scala 117:145]
  assign _T_442 = _T_379 & _T_441; // @[PMP.scala 117:88]
  assign _T_458 = _T_239 & _T_87; // @[PMP.scala 118:113]
  assign _T_459 = _T_458 != 3'h0; // @[PMP.scala 118:146]
  assign _T_460 = _T_232 & _T_459; // @[PMP.scala 118:83]
  assign _T_461 = _T_442 | _T_460; // @[PMP.scala 119:46]
  assign _T_465 = ~_T_39[2:0] & ~io_pmp_5_mask[2:0]; // @[PMP.scala 120:32]
  assign _T_466 = _T_465 == 3'h0; // @[PMP.scala 120:57]
  assign _T_468 = io_pmp_5_cfg_a[1] ? _T_466 : ~_T_461; // @[PMP.scala 121:8]
  assign _T_471 = _T_468 & io_pmp_5_cfg_r; // @[PMP.scala 160:27]
  assign _T_472 = _T_471 | _T_420; // @[PMP.scala 160:41]
  assign _T_473 = _T_468 & io_pmp_5_cfg_w; // @[PMP.scala 161:27]
  assign _T_474 = _T_473 | _T_420; // @[PMP.scala 161:41]
  assign _T_475 = _T_468 & io_pmp_5_cfg_x; // @[PMP.scala 162:27]
  assign _T_476 = _T_475 | _T_420; // @[PMP.scala 162:41]
  assign _T_477_cfg_x = _T_418 ? _T_476 : _T_330_cfg_x; // @[PMP.scala 163:8]
  assign _T_477_cfg_w = _T_418 ? _T_474 : _T_330_cfg_w; // @[PMP.scala 163:8]
  assign _T_477_cfg_r = _T_418 ? _T_472 : _T_330_cfg_r; // @[PMP.scala 163:8]
  assign _T_483 = io_pmp_4_mask | _GEN_0; // @[PMP.scala 62:26]
  assign _T_493 = _T_378 & ~io_pmp_4_mask[31:3]; // @[PMP.scala 57:52]
  assign _T_494 = _T_493 == 29'h0; // @[PMP.scala 57:58]
  assign _T_502 = io_addr[2:0] ^ _T_386; // @[PMP.scala 57:47]
  assign _T_504 = _T_502 & ~_T_483[2:0]; // @[PMP.scala 57:52]
  assign _T_505 = _T_504 == 3'h0; // @[PMP.scala 57:58]
  assign _T_506 = _T_494 & _T_505; // @[PMP.scala 65:16]
  assign _T_513 = {io_pmp_3_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_515 = ~_T_513 | 32'h3; // @[PMP.scala 54:48]
  assign _T_517 = ~_T_515[31:3]; // @[PMP.scala 74:52]
  assign _T_518 = io_addr[31:3] < _T_517; // @[PMP.scala 74:39]
  assign _T_525 = io_addr[31:3] ^ _T_517; // @[PMP.scala 75:41]
  assign _T_526 = _T_525 == 29'h0; // @[PMP.scala 75:69]
  assign _T_533 = ~_T_515[2:0]; // @[PMP.scala 76:64]
  assign _T_534 = _T_87 < _T_533; // @[PMP.scala 76:53]
  assign _T_535 = _T_526 & _T_534; // @[PMP.scala 77:30]
  assign _T_536 = _T_518 | _T_535; // @[PMP.scala 77:16]
  assign _T_560 = io_addr[2:0] < _T_386; // @[PMP.scala 76:53]
  assign _T_561 = _T_379 & _T_560; // @[PMP.scala 77:30]
  assign _T_562 = _T_371 | _T_561; // @[PMP.scala 77:16]
  assign _T_563 = ~_T_536 & _T_562; // @[PMP.scala 88:48]
  assign _T_564 = io_pmp_4_cfg_a[0] & _T_563; // @[PMP.scala 126:61]
  assign _T_565 = io_pmp_4_cfg_a[1] ? _T_506 : _T_564; // @[PMP.scala 126:8]
  assign _T_567 = default_ & ~io_pmp_4_cfg_l; // @[PMP.scala 157:26]
  assign _T_587 = _T_533 & ~io_addr[2:0]; // @[PMP.scala 117:123]
  assign _T_588 = _T_587 != 3'h0; // @[PMP.scala 117:145]
  assign _T_589 = _T_526 & _T_588; // @[PMP.scala 117:88]
  assign _T_605 = _T_386 & _T_87; // @[PMP.scala 118:113]
  assign _T_606 = _T_605 != 3'h0; // @[PMP.scala 118:146]
  assign _T_607 = _T_379 & _T_606; // @[PMP.scala 118:83]
  assign _T_608 = _T_589 | _T_607; // @[PMP.scala 119:46]
  assign _T_612 = ~_T_39[2:0] & ~io_pmp_4_mask[2:0]; // @[PMP.scala 120:32]
  assign _T_613 = _T_612 == 3'h0; // @[PMP.scala 120:57]
  assign _T_615 = io_pmp_4_cfg_a[1] ? _T_613 : ~_T_608; // @[PMP.scala 121:8]
  assign _T_618 = _T_615 & io_pmp_4_cfg_r; // @[PMP.scala 160:27]
  assign _T_619 = _T_618 | _T_567; // @[PMP.scala 160:41]
  assign _T_620 = _T_615 & io_pmp_4_cfg_w; // @[PMP.scala 161:27]
  assign _T_621 = _T_620 | _T_567; // @[PMP.scala 161:41]
  assign _T_622 = _T_615 & io_pmp_4_cfg_x; // @[PMP.scala 162:27]
  assign _T_623 = _T_622 | _T_567; // @[PMP.scala 162:41]
  assign _T_624_cfg_x = _T_565 ? _T_623 : _T_477_cfg_x; // @[PMP.scala 163:8]
  assign _T_624_cfg_w = _T_565 ? _T_621 : _T_477_cfg_w; // @[PMP.scala 163:8]
  assign _T_624_cfg_r = _T_565 ? _T_619 : _T_477_cfg_r; // @[PMP.scala 163:8]
  assign _T_630 = io_pmp_3_mask | _GEN_0; // @[PMP.scala 62:26]
  assign _T_640 = _T_525 & ~io_pmp_3_mask[31:3]; // @[PMP.scala 57:52]
  assign _T_641 = _T_640 == 29'h0; // @[PMP.scala 57:58]
  assign _T_649 = io_addr[2:0] ^ _T_533; // @[PMP.scala 57:47]
  assign _T_651 = _T_649 & ~_T_630[2:0]; // @[PMP.scala 57:52]
  assign _T_652 = _T_651 == 3'h0; // @[PMP.scala 57:58]
  assign _T_653 = _T_641 & _T_652; // @[PMP.scala 65:16]
  assign _T_660 = {io_pmp_2_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_662 = ~_T_660 | 32'h3; // @[PMP.scala 54:48]
  assign _T_664 = ~_T_662[31:3]; // @[PMP.scala 74:52]
  assign _T_665 = io_addr[31:3] < _T_664; // @[PMP.scala 74:39]
  assign _T_672 = io_addr[31:3] ^ _T_664; // @[PMP.scala 75:41]
  assign _T_673 = _T_672 == 29'h0; // @[PMP.scala 75:69]
  assign _T_680 = ~_T_662[2:0]; // @[PMP.scala 76:64]
  assign _T_681 = _T_87 < _T_680; // @[PMP.scala 76:53]
  assign _T_682 = _T_673 & _T_681; // @[PMP.scala 77:30]
  assign _T_683 = _T_665 | _T_682; // @[PMP.scala 77:16]
  assign _T_707 = io_addr[2:0] < _T_533; // @[PMP.scala 76:53]
  assign _T_708 = _T_526 & _T_707; // @[PMP.scala 77:30]
  assign _T_709 = _T_518 | _T_708; // @[PMP.scala 77:16]
  assign _T_710 = ~_T_683 & _T_709; // @[PMP.scala 88:48]
  assign _T_711 = io_pmp_3_cfg_a[0] & _T_710; // @[PMP.scala 126:61]
  assign _T_712 = io_pmp_3_cfg_a[1] ? _T_653 : _T_711; // @[PMP.scala 126:8]
  assign _T_714 = default_ & ~io_pmp_3_cfg_l; // @[PMP.scala 157:26]
  assign _T_734 = _T_680 & ~io_addr[2:0]; // @[PMP.scala 117:123]
  assign _T_735 = _T_734 != 3'h0; // @[PMP.scala 117:145]
  assign _T_736 = _T_673 & _T_735; // @[PMP.scala 117:88]
  assign _T_752 = _T_533 & _T_87; // @[PMP.scala 118:113]
  assign _T_753 = _T_752 != 3'h0; // @[PMP.scala 118:146]
  assign _T_754 = _T_526 & _T_753; // @[PMP.scala 118:83]
  assign _T_755 = _T_736 | _T_754; // @[PMP.scala 119:46]
  assign _T_759 = ~_T_39[2:0] & ~io_pmp_3_mask[2:0]; // @[PMP.scala 120:32]
  assign _T_760 = _T_759 == 3'h0; // @[PMP.scala 120:57]
  assign _T_762 = io_pmp_3_cfg_a[1] ? _T_760 : ~_T_755; // @[PMP.scala 121:8]
  assign _T_765 = _T_762 & io_pmp_3_cfg_r; // @[PMP.scala 160:27]
  assign _T_766 = _T_765 | _T_714; // @[PMP.scala 160:41]
  assign _T_767 = _T_762 & io_pmp_3_cfg_w; // @[PMP.scala 161:27]
  assign _T_768 = _T_767 | _T_714; // @[PMP.scala 161:41]
  assign _T_769 = _T_762 & io_pmp_3_cfg_x; // @[PMP.scala 162:27]
  assign _T_770 = _T_769 | _T_714; // @[PMP.scala 162:41]
  assign _T_771_cfg_x = _T_712 ? _T_770 : _T_624_cfg_x; // @[PMP.scala 163:8]
  assign _T_771_cfg_w = _T_712 ? _T_768 : _T_624_cfg_w; // @[PMP.scala 163:8]
  assign _T_771_cfg_r = _T_712 ? _T_766 : _T_624_cfg_r; // @[PMP.scala 163:8]
  assign _T_777 = io_pmp_2_mask | _GEN_0; // @[PMP.scala 62:26]
  assign _T_787 = _T_672 & ~io_pmp_2_mask[31:3]; // @[PMP.scala 57:52]
  assign _T_788 = _T_787 == 29'h0; // @[PMP.scala 57:58]
  assign _T_796 = io_addr[2:0] ^ _T_680; // @[PMP.scala 57:47]
  assign _T_798 = _T_796 & ~_T_777[2:0]; // @[PMP.scala 57:52]
  assign _T_799 = _T_798 == 3'h0; // @[PMP.scala 57:58]
  assign _T_800 = _T_788 & _T_799; // @[PMP.scala 65:16]
  assign _T_807 = {io_pmp_1_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_809 = ~_T_807 | 32'h3; // @[PMP.scala 54:48]
  assign _T_811 = ~_T_809[31:3]; // @[PMP.scala 74:52]
  assign _T_812 = io_addr[31:3] < _T_811; // @[PMP.scala 74:39]
  assign _T_819 = io_addr[31:3] ^ _T_811; // @[PMP.scala 75:41]
  assign _T_820 = _T_819 == 29'h0; // @[PMP.scala 75:69]
  assign _T_827 = ~_T_809[2:0]; // @[PMP.scala 76:64]
  assign _T_828 = _T_87 < _T_827; // @[PMP.scala 76:53]
  assign _T_829 = _T_820 & _T_828; // @[PMP.scala 77:30]
  assign _T_830 = _T_812 | _T_829; // @[PMP.scala 77:16]
  assign _T_854 = io_addr[2:0] < _T_680; // @[PMP.scala 76:53]
  assign _T_855 = _T_673 & _T_854; // @[PMP.scala 77:30]
  assign _T_856 = _T_665 | _T_855; // @[PMP.scala 77:16]
  assign _T_857 = ~_T_830 & _T_856; // @[PMP.scala 88:48]
  assign _T_858 = io_pmp_2_cfg_a[0] & _T_857; // @[PMP.scala 126:61]
  assign _T_859 = io_pmp_2_cfg_a[1] ? _T_800 : _T_858; // @[PMP.scala 126:8]
  assign _T_861 = default_ & ~io_pmp_2_cfg_l; // @[PMP.scala 157:26]
  assign _T_881 = _T_827 & ~io_addr[2:0]; // @[PMP.scala 117:123]
  assign _T_882 = _T_881 != 3'h0; // @[PMP.scala 117:145]
  assign _T_883 = _T_820 & _T_882; // @[PMP.scala 117:88]
  assign _T_899 = _T_680 & _T_87; // @[PMP.scala 118:113]
  assign _T_900 = _T_899 != 3'h0; // @[PMP.scala 118:146]
  assign _T_901 = _T_673 & _T_900; // @[PMP.scala 118:83]
  assign _T_902 = _T_883 | _T_901; // @[PMP.scala 119:46]
  assign _T_906 = ~_T_39[2:0] & ~io_pmp_2_mask[2:0]; // @[PMP.scala 120:32]
  assign _T_907 = _T_906 == 3'h0; // @[PMP.scala 120:57]
  assign _T_909 = io_pmp_2_cfg_a[1] ? _T_907 : ~_T_902; // @[PMP.scala 121:8]
  assign _T_912 = _T_909 & io_pmp_2_cfg_r; // @[PMP.scala 160:27]
  assign _T_913 = _T_912 | _T_861; // @[PMP.scala 160:41]
  assign _T_914 = _T_909 & io_pmp_2_cfg_w; // @[PMP.scala 161:27]
  assign _T_915 = _T_914 | _T_861; // @[PMP.scala 161:41]
  assign _T_916 = _T_909 & io_pmp_2_cfg_x; // @[PMP.scala 162:27]
  assign _T_917 = _T_916 | _T_861; // @[PMP.scala 162:41]
  assign _T_918_cfg_x = _T_859 ? _T_917 : _T_771_cfg_x; // @[PMP.scala 163:8]
  assign _T_918_cfg_w = _T_859 ? _T_915 : _T_771_cfg_w; // @[PMP.scala 163:8]
  assign _T_918_cfg_r = _T_859 ? _T_913 : _T_771_cfg_r; // @[PMP.scala 163:8]
  assign _T_924 = io_pmp_1_mask | _GEN_0; // @[PMP.scala 62:26]
  assign _T_934 = _T_819 & ~io_pmp_1_mask[31:3]; // @[PMP.scala 57:52]
  assign _T_935 = _T_934 == 29'h0; // @[PMP.scala 57:58]
  assign _T_943 = io_addr[2:0] ^ _T_827; // @[PMP.scala 57:47]
  assign _T_945 = _T_943 & ~_T_924[2:0]; // @[PMP.scala 57:52]
  assign _T_946 = _T_945 == 3'h0; // @[PMP.scala 57:58]
  assign _T_947 = _T_935 & _T_946; // @[PMP.scala 65:16]
  assign _T_954 = {io_pmp_0_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_956 = ~_T_954 | 32'h3; // @[PMP.scala 54:48]
  assign _T_958 = ~_T_956[31:3]; // @[PMP.scala 74:52]
  assign _T_959 = io_addr[31:3] < _T_958; // @[PMP.scala 74:39]
  assign _T_966 = io_addr[31:3] ^ _T_958; // @[PMP.scala 75:41]
  assign _T_967 = _T_966 == 29'h0; // @[PMP.scala 75:69]
  assign _T_974 = ~_T_956[2:0]; // @[PMP.scala 76:64]
  assign _T_975 = _T_87 < _T_974; // @[PMP.scala 76:53]
  assign _T_976 = _T_967 & _T_975; // @[PMP.scala 77:30]
  assign _T_977 = _T_959 | _T_976; // @[PMP.scala 77:16]
  assign _T_1001 = io_addr[2:0] < _T_827; // @[PMP.scala 76:53]
  assign _T_1002 = _T_820 & _T_1001; // @[PMP.scala 77:30]
  assign _T_1003 = _T_812 | _T_1002; // @[PMP.scala 77:16]
  assign _T_1004 = ~_T_977 & _T_1003; // @[PMP.scala 88:48]
  assign _T_1005 = io_pmp_1_cfg_a[0] & _T_1004; // @[PMP.scala 126:61]
  assign _T_1006 = io_pmp_1_cfg_a[1] ? _T_947 : _T_1005; // @[PMP.scala 126:8]
  assign _T_1008 = default_ & ~io_pmp_1_cfg_l; // @[PMP.scala 157:26]
  assign _T_1028 = _T_974 & ~io_addr[2:0]; // @[PMP.scala 117:123]
  assign _T_1029 = _T_1028 != 3'h0; // @[PMP.scala 117:145]
  assign _T_1030 = _T_967 & _T_1029; // @[PMP.scala 117:88]
  assign _T_1046 = _T_827 & _T_87; // @[PMP.scala 118:113]
  assign _T_1047 = _T_1046 != 3'h0; // @[PMP.scala 118:146]
  assign _T_1048 = _T_820 & _T_1047; // @[PMP.scala 118:83]
  assign _T_1049 = _T_1030 | _T_1048; // @[PMP.scala 119:46]
  assign _T_1053 = ~_T_39[2:0] & ~io_pmp_1_mask[2:0]; // @[PMP.scala 120:32]
  assign _T_1054 = _T_1053 == 3'h0; // @[PMP.scala 120:57]
  assign _T_1056 = io_pmp_1_cfg_a[1] ? _T_1054 : ~_T_1049; // @[PMP.scala 121:8]
  assign _T_1059 = _T_1056 & io_pmp_1_cfg_r; // @[PMP.scala 160:27]
  assign _T_1060 = _T_1059 | _T_1008; // @[PMP.scala 160:41]
  assign _T_1061 = _T_1056 & io_pmp_1_cfg_w; // @[PMP.scala 161:27]
  assign _T_1062 = _T_1061 | _T_1008; // @[PMP.scala 161:41]
  assign _T_1063 = _T_1056 & io_pmp_1_cfg_x; // @[PMP.scala 162:27]
  assign _T_1064 = _T_1063 | _T_1008; // @[PMP.scala 162:41]
  assign _T_1065_cfg_x = _T_1006 ? _T_1064 : _T_918_cfg_x; // @[PMP.scala 163:8]
  assign _T_1065_cfg_w = _T_1006 ? _T_1062 : _T_918_cfg_w; // @[PMP.scala 163:8]
  assign _T_1065_cfg_r = _T_1006 ? _T_1060 : _T_918_cfg_r; // @[PMP.scala 163:8]
  assign _T_1071 = io_pmp_0_mask | _GEN_0; // @[PMP.scala 62:26]
  assign _T_1081 = _T_966 & ~io_pmp_0_mask[31:3]; // @[PMP.scala 57:52]
  assign _T_1082 = _T_1081 == 29'h0; // @[PMP.scala 57:58]
  assign _T_1090 = io_addr[2:0] ^ _T_974; // @[PMP.scala 57:47]
  assign _T_1092 = _T_1090 & ~_T_1071[2:0]; // @[PMP.scala 57:52]
  assign _T_1093 = _T_1092 == 3'h0; // @[PMP.scala 57:58]
  assign _T_1094 = _T_1082 & _T_1093; // @[PMP.scala 65:16]
  assign _T_1148 = io_addr[2:0] < _T_974; // @[PMP.scala 76:53]
  assign _T_1149 = _T_967 & _T_1148; // @[PMP.scala 77:30]
  assign _T_1150 = _T_959 | _T_1149; // @[PMP.scala 77:16]
  assign _T_1152 = io_pmp_0_cfg_a[0] & _T_1150; // @[PMP.scala 126:61]
  assign _T_1153 = io_pmp_0_cfg_a[1] ? _T_1094 : _T_1152; // @[PMP.scala 126:8]
  assign _T_1155 = default_ & ~io_pmp_0_cfg_l; // @[PMP.scala 157:26]
  assign _T_1193 = _T_974 & _T_87; // @[PMP.scala 118:113]
  assign _T_1194 = _T_1193 != 3'h0; // @[PMP.scala 118:146]
  assign _T_1195 = _T_967 & _T_1194; // @[PMP.scala 118:83]
  assign _T_1200 = ~_T_39[2:0] & ~io_pmp_0_mask[2:0]; // @[PMP.scala 120:32]
  assign _T_1201 = _T_1200 == 3'h0; // @[PMP.scala 120:57]
  assign _T_1203 = io_pmp_0_cfg_a[1] ? _T_1201 : ~_T_1195; // @[PMP.scala 121:8]
  assign _T_1206 = _T_1203 & io_pmp_0_cfg_r; // @[PMP.scala 160:27]
  assign _T_1207 = _T_1206 | _T_1155; // @[PMP.scala 160:41]
  assign _T_1208 = _T_1203 & io_pmp_0_cfg_w; // @[PMP.scala 161:27]
  assign _T_1209 = _T_1208 | _T_1155; // @[PMP.scala 161:41]
  assign _T_1210 = _T_1203 & io_pmp_0_cfg_x; // @[PMP.scala 162:27]
  assign _T_1211 = _T_1210 | _T_1155; // @[PMP.scala 162:41]
  assign io_r = _T_1153 ? _T_1207 : _T_1065_cfg_r; // @[PMP.scala 166:8]
  assign io_w = _T_1153 ? _T_1209 : _T_1065_cfg_w; // @[PMP.scala 167:8]
  assign io_x = _T_1153 ? _T_1211 : _T_1065_cfg_x; // @[PMP.scala 168:8]
  assign PMPChecker_covSum = 30'h0;
  assign io_covSum = PMPChecker_covSum;
  assign metaAssert = 1'h0;
endmodule
module PMPChecker_1(
  input  [1:0]  io_prv,
  input         io_pmp_0_cfg_l,
  input  [1:0]  io_pmp_0_cfg_a,
  input         io_pmp_0_cfg_x,
  input         io_pmp_0_cfg_w,
  input         io_pmp_0_cfg_r,
  input  [29:0] io_pmp_0_addr,
  input  [31:0] io_pmp_0_mask,
  input         io_pmp_1_cfg_l,
  input  [1:0]  io_pmp_1_cfg_a,
  input         io_pmp_1_cfg_x,
  input         io_pmp_1_cfg_w,
  input         io_pmp_1_cfg_r,
  input  [29:0] io_pmp_1_addr,
  input  [31:0] io_pmp_1_mask,
  input         io_pmp_2_cfg_l,
  input  [1:0]  io_pmp_2_cfg_a,
  input         io_pmp_2_cfg_x,
  input         io_pmp_2_cfg_w,
  input         io_pmp_2_cfg_r,
  input  [29:0] io_pmp_2_addr,
  input  [31:0] io_pmp_2_mask,
  input         io_pmp_3_cfg_l,
  input  [1:0]  io_pmp_3_cfg_a,
  input         io_pmp_3_cfg_x,
  input         io_pmp_3_cfg_w,
  input         io_pmp_3_cfg_r,
  input  [29:0] io_pmp_3_addr,
  input  [31:0] io_pmp_3_mask,
  input         io_pmp_4_cfg_l,
  input  [1:0]  io_pmp_4_cfg_a,
  input         io_pmp_4_cfg_x,
  input         io_pmp_4_cfg_w,
  input         io_pmp_4_cfg_r,
  input  [29:0] io_pmp_4_addr,
  input  [31:0] io_pmp_4_mask,
  input         io_pmp_5_cfg_l,
  input  [1:0]  io_pmp_5_cfg_a,
  input         io_pmp_5_cfg_x,
  input         io_pmp_5_cfg_w,
  input         io_pmp_5_cfg_r,
  input  [29:0] io_pmp_5_addr,
  input  [31:0] io_pmp_5_mask,
  input         io_pmp_6_cfg_l,
  input  [1:0]  io_pmp_6_cfg_a,
  input         io_pmp_6_cfg_x,
  input         io_pmp_6_cfg_w,
  input         io_pmp_6_cfg_r,
  input  [29:0] io_pmp_6_addr,
  input  [31:0] io_pmp_6_mask,
  input         io_pmp_7_cfg_l,
  input  [1:0]  io_pmp_7_cfg_a,
  input         io_pmp_7_cfg_x,
  input         io_pmp_7_cfg_w,
  input         io_pmp_7_cfg_r,
  input  [29:0] io_pmp_7_addr,
  input  [31:0] io_pmp_7_mask,
  input  [31:0] io_addr,
  output        io_r,
  output        io_w,
  output        io_x,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  default_; // @[PMP.scala 149:56]
  wire [31:0] _T_38; // @[PMP.scala 54:36]
  wire [31:0] _T_40; // @[PMP.scala 54:48]
  wire [31:0] _T_42; // @[PMP.scala 57:47]
  wire [31:0] _T_44; // @[PMP.scala 57:52]
  wire  _T_45; // @[PMP.scala 57:58]
  wire [31:0] _T_51; // @[PMP.scala 54:36]
  wire [31:0] _T_53; // @[PMP.scala 54:48]
  wire  _T_55; // @[PMP.scala 71:9]
  wire  _T_61; // @[PMP.scala 71:9]
  wire  _T_62; // @[PMP.scala 88:48]
  wire  _T_63; // @[PMP.scala 126:61]
  wire  _T_64; // @[PMP.scala 126:8]
  wire  _T_66; // @[PMP.scala 157:26]
  wire  _T_70; // @[PMP.scala 160:41]
  wire  _T_72; // @[PMP.scala 161:41]
  wire  _T_74; // @[PMP.scala 162:41]
  wire  _T_75_cfg_x; // @[PMP.scala 163:8]
  wire  _T_75_cfg_w; // @[PMP.scala 163:8]
  wire  _T_75_cfg_r; // @[PMP.scala 163:8]
  wire [31:0] _T_81; // @[PMP.scala 57:47]
  wire [31:0] _T_83; // @[PMP.scala 57:52]
  wire  _T_84; // @[PMP.scala 57:58]
  wire [31:0] _T_90; // @[PMP.scala 54:36]
  wire [31:0] _T_92; // @[PMP.scala 54:48]
  wire  _T_94; // @[PMP.scala 71:9]
  wire  _T_101; // @[PMP.scala 88:48]
  wire  _T_102; // @[PMP.scala 126:61]
  wire  _T_103; // @[PMP.scala 126:8]
  wire  _T_105; // @[PMP.scala 157:26]
  wire  _T_109; // @[PMP.scala 160:41]
  wire  _T_111; // @[PMP.scala 161:41]
  wire  _T_113; // @[PMP.scala 162:41]
  wire  _T_114_cfg_x; // @[PMP.scala 163:8]
  wire  _T_114_cfg_w; // @[PMP.scala 163:8]
  wire  _T_114_cfg_r; // @[PMP.scala 163:8]
  wire [31:0] _T_120; // @[PMP.scala 57:47]
  wire [31:0] _T_122; // @[PMP.scala 57:52]
  wire  _T_123; // @[PMP.scala 57:58]
  wire [31:0] _T_129; // @[PMP.scala 54:36]
  wire [31:0] _T_131; // @[PMP.scala 54:48]
  wire  _T_133; // @[PMP.scala 71:9]
  wire  _T_140; // @[PMP.scala 88:48]
  wire  _T_141; // @[PMP.scala 126:61]
  wire  _T_142; // @[PMP.scala 126:8]
  wire  _T_144; // @[PMP.scala 157:26]
  wire  _T_148; // @[PMP.scala 160:41]
  wire  _T_150; // @[PMP.scala 161:41]
  wire  _T_152; // @[PMP.scala 162:41]
  wire  _T_153_cfg_x; // @[PMP.scala 163:8]
  wire  _T_153_cfg_w; // @[PMP.scala 163:8]
  wire  _T_153_cfg_r; // @[PMP.scala 163:8]
  wire [31:0] _T_159; // @[PMP.scala 57:47]
  wire [31:0] _T_161; // @[PMP.scala 57:52]
  wire  _T_162; // @[PMP.scala 57:58]
  wire [31:0] _T_168; // @[PMP.scala 54:36]
  wire [31:0] _T_170; // @[PMP.scala 54:48]
  wire  _T_172; // @[PMP.scala 71:9]
  wire  _T_179; // @[PMP.scala 88:48]
  wire  _T_180; // @[PMP.scala 126:61]
  wire  _T_181; // @[PMP.scala 126:8]
  wire  _T_183; // @[PMP.scala 157:26]
  wire  _T_187; // @[PMP.scala 160:41]
  wire  _T_189; // @[PMP.scala 161:41]
  wire  _T_191; // @[PMP.scala 162:41]
  wire  _T_192_cfg_x; // @[PMP.scala 163:8]
  wire  _T_192_cfg_w; // @[PMP.scala 163:8]
  wire  _T_192_cfg_r; // @[PMP.scala 163:8]
  wire [31:0] _T_198; // @[PMP.scala 57:47]
  wire [31:0] _T_200; // @[PMP.scala 57:52]
  wire  _T_201; // @[PMP.scala 57:58]
  wire [31:0] _T_207; // @[PMP.scala 54:36]
  wire [31:0] _T_209; // @[PMP.scala 54:48]
  wire  _T_211; // @[PMP.scala 71:9]
  wire  _T_218; // @[PMP.scala 88:48]
  wire  _T_219; // @[PMP.scala 126:61]
  wire  _T_220; // @[PMP.scala 126:8]
  wire  _T_222; // @[PMP.scala 157:26]
  wire  _T_226; // @[PMP.scala 160:41]
  wire  _T_228; // @[PMP.scala 161:41]
  wire  _T_230; // @[PMP.scala 162:41]
  wire  _T_231_cfg_x; // @[PMP.scala 163:8]
  wire  _T_231_cfg_w; // @[PMP.scala 163:8]
  wire  _T_231_cfg_r; // @[PMP.scala 163:8]
  wire [31:0] _T_237; // @[PMP.scala 57:47]
  wire [31:0] _T_239; // @[PMP.scala 57:52]
  wire  _T_240; // @[PMP.scala 57:58]
  wire [31:0] _T_246; // @[PMP.scala 54:36]
  wire [31:0] _T_248; // @[PMP.scala 54:48]
  wire  _T_250; // @[PMP.scala 71:9]
  wire  _T_257; // @[PMP.scala 88:48]
  wire  _T_258; // @[PMP.scala 126:61]
  wire  _T_259; // @[PMP.scala 126:8]
  wire  _T_261; // @[PMP.scala 157:26]
  wire  _T_265; // @[PMP.scala 160:41]
  wire  _T_267; // @[PMP.scala 161:41]
  wire  _T_269; // @[PMP.scala 162:41]
  wire  _T_270_cfg_x; // @[PMP.scala 163:8]
  wire  _T_270_cfg_w; // @[PMP.scala 163:8]
  wire  _T_270_cfg_r; // @[PMP.scala 163:8]
  wire [31:0] _T_276; // @[PMP.scala 57:47]
  wire [31:0] _T_278; // @[PMP.scala 57:52]
  wire  _T_279; // @[PMP.scala 57:58]
  wire [31:0] _T_285; // @[PMP.scala 54:36]
  wire [31:0] _T_287; // @[PMP.scala 54:48]
  wire  _T_289; // @[PMP.scala 71:9]
  wire  _T_296; // @[PMP.scala 88:48]
  wire  _T_297; // @[PMP.scala 126:61]
  wire  _T_298; // @[PMP.scala 126:8]
  wire  _T_300; // @[PMP.scala 157:26]
  wire  _T_304; // @[PMP.scala 160:41]
  wire  _T_306; // @[PMP.scala 161:41]
  wire  _T_308; // @[PMP.scala 162:41]
  wire  _T_309_cfg_x; // @[PMP.scala 163:8]
  wire  _T_309_cfg_w; // @[PMP.scala 163:8]
  wire  _T_309_cfg_r; // @[PMP.scala 163:8]
  wire [31:0] _T_315; // @[PMP.scala 57:47]
  wire [31:0] _T_317; // @[PMP.scala 57:52]
  wire  _T_318; // @[PMP.scala 57:58]
  wire  _T_336; // @[PMP.scala 126:61]
  wire  _T_337; // @[PMP.scala 126:8]
  wire  _T_339; // @[PMP.scala 157:26]
  wire  _T_343; // @[PMP.scala 160:41]
  wire  _T_345; // @[PMP.scala 161:41]
  wire  _T_347; // @[PMP.scala 162:41]
  wire [29:0] PMPChecker_1_covSum;
  assign default_ = io_prv > 2'h1; // @[PMP.scala 149:56]
  assign _T_38 = {io_pmp_7_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_40 = ~_T_38 | 32'h3; // @[PMP.scala 54:48]
  assign _T_42 = io_addr ^ ~_T_40; // @[PMP.scala 57:47]
  assign _T_44 = _T_42 & ~io_pmp_7_mask; // @[PMP.scala 57:52]
  assign _T_45 = _T_44 == 32'h0; // @[PMP.scala 57:58]
  assign _T_51 = {io_pmp_6_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_53 = ~_T_51 | 32'h3; // @[PMP.scala 54:48]
  assign _T_55 = io_addr < ~_T_53; // @[PMP.scala 71:9]
  assign _T_61 = io_addr < ~_T_40; // @[PMP.scala 71:9]
  assign _T_62 = ~_T_55 & _T_61; // @[PMP.scala 88:48]
  assign _T_63 = io_pmp_7_cfg_a[0] & _T_62; // @[PMP.scala 126:61]
  assign _T_64 = io_pmp_7_cfg_a[1] ? _T_45 : _T_63; // @[PMP.scala 126:8]
  assign _T_66 = default_ & ~io_pmp_7_cfg_l; // @[PMP.scala 157:26]
  assign _T_70 = io_pmp_7_cfg_r | _T_66; // @[PMP.scala 160:41]
  assign _T_72 = io_pmp_7_cfg_w | _T_66; // @[PMP.scala 161:41]
  assign _T_74 = io_pmp_7_cfg_x | _T_66; // @[PMP.scala 162:41]
  assign _T_75_cfg_x = _T_64 ? _T_74 : default_; // @[PMP.scala 163:8]
  assign _T_75_cfg_w = _T_64 ? _T_72 : default_; // @[PMP.scala 163:8]
  assign _T_75_cfg_r = _T_64 ? _T_70 : default_; // @[PMP.scala 163:8]
  assign _T_81 = io_addr ^ ~_T_53; // @[PMP.scala 57:47]
  assign _T_83 = _T_81 & ~io_pmp_6_mask; // @[PMP.scala 57:52]
  assign _T_84 = _T_83 == 32'h0; // @[PMP.scala 57:58]
  assign _T_90 = {io_pmp_5_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_92 = ~_T_90 | 32'h3; // @[PMP.scala 54:48]
  assign _T_94 = io_addr < ~_T_92; // @[PMP.scala 71:9]
  assign _T_101 = ~_T_94 & _T_55; // @[PMP.scala 88:48]
  assign _T_102 = io_pmp_6_cfg_a[0] & _T_101; // @[PMP.scala 126:61]
  assign _T_103 = io_pmp_6_cfg_a[1] ? _T_84 : _T_102; // @[PMP.scala 126:8]
  assign _T_105 = default_ & ~io_pmp_6_cfg_l; // @[PMP.scala 157:26]
  assign _T_109 = io_pmp_6_cfg_r | _T_105; // @[PMP.scala 160:41]
  assign _T_111 = io_pmp_6_cfg_w | _T_105; // @[PMP.scala 161:41]
  assign _T_113 = io_pmp_6_cfg_x | _T_105; // @[PMP.scala 162:41]
  assign _T_114_cfg_x = _T_103 ? _T_113 : _T_75_cfg_x; // @[PMP.scala 163:8]
  assign _T_114_cfg_w = _T_103 ? _T_111 : _T_75_cfg_w; // @[PMP.scala 163:8]
  assign _T_114_cfg_r = _T_103 ? _T_109 : _T_75_cfg_r; // @[PMP.scala 163:8]
  assign _T_120 = io_addr ^ ~_T_92; // @[PMP.scala 57:47]
  assign _T_122 = _T_120 & ~io_pmp_5_mask; // @[PMP.scala 57:52]
  assign _T_123 = _T_122 == 32'h0; // @[PMP.scala 57:58]
  assign _T_129 = {io_pmp_4_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_131 = ~_T_129 | 32'h3; // @[PMP.scala 54:48]
  assign _T_133 = io_addr < ~_T_131; // @[PMP.scala 71:9]
  assign _T_140 = ~_T_133 & _T_94; // @[PMP.scala 88:48]
  assign _T_141 = io_pmp_5_cfg_a[0] & _T_140; // @[PMP.scala 126:61]
  assign _T_142 = io_pmp_5_cfg_a[1] ? _T_123 : _T_141; // @[PMP.scala 126:8]
  assign _T_144 = default_ & ~io_pmp_5_cfg_l; // @[PMP.scala 157:26]
  assign _T_148 = io_pmp_5_cfg_r | _T_144; // @[PMP.scala 160:41]
  assign _T_150 = io_pmp_5_cfg_w | _T_144; // @[PMP.scala 161:41]
  assign _T_152 = io_pmp_5_cfg_x | _T_144; // @[PMP.scala 162:41]
  assign _T_153_cfg_x = _T_142 ? _T_152 : _T_114_cfg_x; // @[PMP.scala 163:8]
  assign _T_153_cfg_w = _T_142 ? _T_150 : _T_114_cfg_w; // @[PMP.scala 163:8]
  assign _T_153_cfg_r = _T_142 ? _T_148 : _T_114_cfg_r; // @[PMP.scala 163:8]
  assign _T_159 = io_addr ^ ~_T_131; // @[PMP.scala 57:47]
  assign _T_161 = _T_159 & ~io_pmp_4_mask; // @[PMP.scala 57:52]
  assign _T_162 = _T_161 == 32'h0; // @[PMP.scala 57:58]
  assign _T_168 = {io_pmp_3_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_170 = ~_T_168 | 32'h3; // @[PMP.scala 54:48]
  assign _T_172 = io_addr < ~_T_170; // @[PMP.scala 71:9]
  assign _T_179 = ~_T_172 & _T_133; // @[PMP.scala 88:48]
  assign _T_180 = io_pmp_4_cfg_a[0] & _T_179; // @[PMP.scala 126:61]
  assign _T_181 = io_pmp_4_cfg_a[1] ? _T_162 : _T_180; // @[PMP.scala 126:8]
  assign _T_183 = default_ & ~io_pmp_4_cfg_l; // @[PMP.scala 157:26]
  assign _T_187 = io_pmp_4_cfg_r | _T_183; // @[PMP.scala 160:41]
  assign _T_189 = io_pmp_4_cfg_w | _T_183; // @[PMP.scala 161:41]
  assign _T_191 = io_pmp_4_cfg_x | _T_183; // @[PMP.scala 162:41]
  assign _T_192_cfg_x = _T_181 ? _T_191 : _T_153_cfg_x; // @[PMP.scala 163:8]
  assign _T_192_cfg_w = _T_181 ? _T_189 : _T_153_cfg_w; // @[PMP.scala 163:8]
  assign _T_192_cfg_r = _T_181 ? _T_187 : _T_153_cfg_r; // @[PMP.scala 163:8]
  assign _T_198 = io_addr ^ ~_T_170; // @[PMP.scala 57:47]
  assign _T_200 = _T_198 & ~io_pmp_3_mask; // @[PMP.scala 57:52]
  assign _T_201 = _T_200 == 32'h0; // @[PMP.scala 57:58]
  assign _T_207 = {io_pmp_2_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_209 = ~_T_207 | 32'h3; // @[PMP.scala 54:48]
  assign _T_211 = io_addr < ~_T_209; // @[PMP.scala 71:9]
  assign _T_218 = ~_T_211 & _T_172; // @[PMP.scala 88:48]
  assign _T_219 = io_pmp_3_cfg_a[0] & _T_218; // @[PMP.scala 126:61]
  assign _T_220 = io_pmp_3_cfg_a[1] ? _T_201 : _T_219; // @[PMP.scala 126:8]
  assign _T_222 = default_ & ~io_pmp_3_cfg_l; // @[PMP.scala 157:26]
  assign _T_226 = io_pmp_3_cfg_r | _T_222; // @[PMP.scala 160:41]
  assign _T_228 = io_pmp_3_cfg_w | _T_222; // @[PMP.scala 161:41]
  assign _T_230 = io_pmp_3_cfg_x | _T_222; // @[PMP.scala 162:41]
  assign _T_231_cfg_x = _T_220 ? _T_230 : _T_192_cfg_x; // @[PMP.scala 163:8]
  assign _T_231_cfg_w = _T_220 ? _T_228 : _T_192_cfg_w; // @[PMP.scala 163:8]
  assign _T_231_cfg_r = _T_220 ? _T_226 : _T_192_cfg_r; // @[PMP.scala 163:8]
  assign _T_237 = io_addr ^ ~_T_209; // @[PMP.scala 57:47]
  assign _T_239 = _T_237 & ~io_pmp_2_mask; // @[PMP.scala 57:52]
  assign _T_240 = _T_239 == 32'h0; // @[PMP.scala 57:58]
  assign _T_246 = {io_pmp_1_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_248 = ~_T_246 | 32'h3; // @[PMP.scala 54:48]
  assign _T_250 = io_addr < ~_T_248; // @[PMP.scala 71:9]
  assign _T_257 = ~_T_250 & _T_211; // @[PMP.scala 88:48]
  assign _T_258 = io_pmp_2_cfg_a[0] & _T_257; // @[PMP.scala 126:61]
  assign _T_259 = io_pmp_2_cfg_a[1] ? _T_240 : _T_258; // @[PMP.scala 126:8]
  assign _T_261 = default_ & ~io_pmp_2_cfg_l; // @[PMP.scala 157:26]
  assign _T_265 = io_pmp_2_cfg_r | _T_261; // @[PMP.scala 160:41]
  assign _T_267 = io_pmp_2_cfg_w | _T_261; // @[PMP.scala 161:41]
  assign _T_269 = io_pmp_2_cfg_x | _T_261; // @[PMP.scala 162:41]
  assign _T_270_cfg_x = _T_259 ? _T_269 : _T_231_cfg_x; // @[PMP.scala 163:8]
  assign _T_270_cfg_w = _T_259 ? _T_267 : _T_231_cfg_w; // @[PMP.scala 163:8]
  assign _T_270_cfg_r = _T_259 ? _T_265 : _T_231_cfg_r; // @[PMP.scala 163:8]
  assign _T_276 = io_addr ^ ~_T_248; // @[PMP.scala 57:47]
  assign _T_278 = _T_276 & ~io_pmp_1_mask; // @[PMP.scala 57:52]
  assign _T_279 = _T_278 == 32'h0; // @[PMP.scala 57:58]
  assign _T_285 = {io_pmp_0_addr, 2'h0}; // @[PMP.scala 54:36]
  assign _T_287 = ~_T_285 | 32'h3; // @[PMP.scala 54:48]
  assign _T_289 = io_addr < ~_T_287; // @[PMP.scala 71:9]
  assign _T_296 = ~_T_289 & _T_250; // @[PMP.scala 88:48]
  assign _T_297 = io_pmp_1_cfg_a[0] & _T_296; // @[PMP.scala 126:61]
  assign _T_298 = io_pmp_1_cfg_a[1] ? _T_279 : _T_297; // @[PMP.scala 126:8]
  assign _T_300 = default_ & ~io_pmp_1_cfg_l; // @[PMP.scala 157:26]
  assign _T_304 = io_pmp_1_cfg_r | _T_300; // @[PMP.scala 160:41]
  assign _T_306 = io_pmp_1_cfg_w | _T_300; // @[PMP.scala 161:41]
  assign _T_308 = io_pmp_1_cfg_x | _T_300; // @[PMP.scala 162:41]
  assign _T_309_cfg_x = _T_298 ? _T_308 : _T_270_cfg_x; // @[PMP.scala 163:8]
  assign _T_309_cfg_w = _T_298 ? _T_306 : _T_270_cfg_w; // @[PMP.scala 163:8]
  assign _T_309_cfg_r = _T_298 ? _T_304 : _T_270_cfg_r; // @[PMP.scala 163:8]
  assign _T_315 = io_addr ^ ~_T_287; // @[PMP.scala 57:47]
  assign _T_317 = _T_315 & ~io_pmp_0_mask; // @[PMP.scala 57:52]
  assign _T_318 = _T_317 == 32'h0; // @[PMP.scala 57:58]
  assign _T_336 = io_pmp_0_cfg_a[0] & _T_289; // @[PMP.scala 126:61]
  assign _T_337 = io_pmp_0_cfg_a[1] ? _T_318 : _T_336; // @[PMP.scala 126:8]
  assign _T_339 = default_ & ~io_pmp_0_cfg_l; // @[PMP.scala 157:26]
  assign _T_343 = io_pmp_0_cfg_r | _T_339; // @[PMP.scala 160:41]
  assign _T_345 = io_pmp_0_cfg_w | _T_339; // @[PMP.scala 161:41]
  assign _T_347 = io_pmp_0_cfg_x | _T_339; // @[PMP.scala 162:41]
  assign io_r = _T_337 ? _T_343 : _T_309_cfg_r; // @[PMP.scala 166:8]
  assign io_w = _T_337 ? _T_345 : _T_309_cfg_w; // @[PMP.scala 167:8]
  assign io_x = _T_337 ? _T_347 : _T_309_cfg_x; // @[PMP.scala 168:8]
  assign PMPChecker_1_covSum = 30'h0;
  assign io_covSum = PMPChecker_1_covSum;
  assign metaAssert = 1'h0;
endmodule
module MulAddRecFNPipe(
  input         clock,
  input         reset,
  input         io_validin,
  input  [1:0]  io_op,
  input  [32:0] io_a,
  input  [32:0] io_b,
  input  [32:0] io_c,
  input  [2:0]  io_roundingMode,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [1:0] mulAddRecFNToRaw_preMul_io_op; // @[FPU.scala 580:15]
  wire [32:0] mulAddRecFNToRaw_preMul_io_a; // @[FPU.scala 580:15]
  wire [32:0] mulAddRecFNToRaw_preMul_io_b; // @[FPU.scala 580:15]
  wire [32:0] mulAddRecFNToRaw_preMul_io_c; // @[FPU.scala 580:15]
  wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddA; // @[FPU.scala 580:15]
  wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddB; // @[FPU.scala 580:15]
  wire [47:0] mulAddRecFNToRaw_preMul_io_mulAddC; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[FPU.scala 580:15]
  wire [9:0] mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[FPU.scala 580:15]
  wire [4:0] mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[FPU.scala 580:15]
  wire [25:0] mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[FPU.scala 580:15]
  wire [29:0] mulAddRecFNToRaw_preMul_io_covSum; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_metaAssert; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_signProd; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC; // @[FPU.scala 582:15]
  wire [9:0] mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant; // @[FPU.scala 582:15]
  wire [4:0] mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist; // @[FPU.scala 582:15]
  wire [25:0] mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC; // @[FPU.scala 582:15]
  wire [48:0] mulAddRecFNToRaw_postMul_io_mulAddResult; // @[FPU.scala 582:15]
  wire [2:0] mulAddRecFNToRaw_postMul_io_roundingMode; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_invalidExc; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[FPU.scala 582:15]
  wire [9:0] mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[FPU.scala 582:15]
  wire [26:0] mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[FPU.scala 582:15]
  wire [29:0] mulAddRecFNToRaw_postMul_io_covSum; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_metaAssert; // @[FPU.scala 582:15]
  wire  roundRawFNToRecFN_io_invalidExc; // @[FPU.scala 608:35]
  wire  roundRawFNToRecFN_io_infiniteExc; // @[FPU.scala 608:35]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[FPU.scala 608:35]
  wire  roundRawFNToRecFN_io_in_isInf; // @[FPU.scala 608:35]
  wire  roundRawFNToRecFN_io_in_isZero; // @[FPU.scala 608:35]
  wire  roundRawFNToRecFN_io_in_sign; // @[FPU.scala 608:35]
  wire [9:0] roundRawFNToRecFN_io_in_sExp; // @[FPU.scala 608:35]
  wire [26:0] roundRawFNToRecFN_io_in_sig; // @[FPU.scala 608:35]
  wire [2:0] roundRawFNToRecFN_io_roundingMode; // @[FPU.scala 608:35]
  wire  roundRawFNToRecFN_io_detectTininess; // @[FPU.scala 608:35]
  wire [32:0] roundRawFNToRecFN_io_out; // @[FPU.scala 608:35]
  wire [4:0] roundRawFNToRecFN_io_exceptionFlags; // @[FPU.scala 608:35]
  wire [29:0] roundRawFNToRecFN_io_covSum; // @[FPU.scala 608:35]
  wire  roundRawFNToRecFN_metaAssert; // @[FPU.scala 608:35]
  wire [47:0] _T_14; // @[FPU.scala 590:45]
  wire [48:0] mulAddResult; // @[FPU.scala 591:50]
  reg  _T_21_isSigNaNAny; // @[Reg.scala 11:16]
  reg [31:0] _RAND_0;
  reg  _T_21_isNaNAOrB; // @[Reg.scala 11:16]
  reg [31:0] _RAND_1;
  reg  _T_21_isInfA; // @[Reg.scala 11:16]
  reg [31:0] _RAND_2;
  reg  _T_21_isZeroA; // @[Reg.scala 11:16]
  reg [31:0] _RAND_3;
  reg  _T_21_isInfB; // @[Reg.scala 11:16]
  reg [31:0] _RAND_4;
  reg  _T_21_isZeroB; // @[Reg.scala 11:16]
  reg [31:0] _RAND_5;
  reg  _T_21_signProd; // @[Reg.scala 11:16]
  reg [31:0] _RAND_6;
  reg  _T_21_isNaNC; // @[Reg.scala 11:16]
  reg [31:0] _RAND_7;
  reg  _T_21_isInfC; // @[Reg.scala 11:16]
  reg [31:0] _RAND_8;
  reg  _T_21_isZeroC; // @[Reg.scala 11:16]
  reg [31:0] _RAND_9;
  reg [9:0] _T_21_sExpSum; // @[Reg.scala 11:16]
  reg [31:0] _RAND_10;
  reg  _T_21_doSubMags; // @[Reg.scala 11:16]
  reg [31:0] _RAND_11;
  reg  _T_21_CIsDominant; // @[Reg.scala 11:16]
  reg [31:0] _RAND_12;
  reg [4:0] _T_21_CDom_CAlignDist; // @[Reg.scala 11:16]
  reg [31:0] _RAND_13;
  reg [25:0] _T_21_highAlignedSigC; // @[Reg.scala 11:16]
  reg [31:0] _RAND_14;
  reg  _T_21_bit0AlignedSigC; // @[Reg.scala 11:16]
  reg [31:0] _RAND_15;
  reg [48:0] _T_30; // @[Reg.scala 11:16]
  reg [63:0] _RAND_16;
  reg [2:0] _T_39; // @[Reg.scala 11:16]
  reg [31:0] _RAND_17;
  reg [2:0] roundingMode_stage0; // @[Reg.scala 11:16]
  reg [31:0] _RAND_18;
  reg  detectTininess_stage0; // @[Reg.scala 11:16]
  reg [31:0] _RAND_19;
  reg  valid_stage0; // @[Valid.scala 48:22]
  reg [31:0] _RAND_20;
  reg  _T_75; // @[Reg.scala 11:16]
  reg [31:0] _RAND_21;
  reg  _T_84_isNaN; // @[Reg.scala 11:16]
  reg [31:0] _RAND_22;
  reg  _T_84_isInf; // @[Reg.scala 11:16]
  reg [31:0] _RAND_23;
  reg  _T_84_isZero; // @[Reg.scala 11:16]
  reg [31:0] _RAND_24;
  reg  _T_84_sign; // @[Reg.scala 11:16]
  reg [31:0] _RAND_25;
  reg [9:0] _T_84_sExp; // @[Reg.scala 11:16]
  reg [31:0] _RAND_26;
  reg [26:0] _T_84_sig; // @[Reg.scala 11:16]
  reg [31:0] _RAND_27;
  reg [2:0] _T_93; // @[Reg.scala 11:16]
  reg [31:0] _RAND_28;
  reg  _T_102; // @[Reg.scala 11:16]
  reg [31:0] _RAND_29;
  reg  MulAddRecFNPipe_state; // @[Register tracking MulAddRecFNPipe state]
  reg [31:0] _RAND_30;
  reg  MulAddRecFNPipe_cov [0:1]; // @[Coverage map for MulAddRecFNPipe]
  reg [31:0] _RAND_31;
  wire  MulAddRecFNPipe_cov_read_data; // @[Coverage map for MulAddRecFNPipe]
  wire  MulAddRecFNPipe_cov_read_addr; // @[Coverage map for MulAddRecFNPipe]
  wire  MulAddRecFNPipe_cov_write_data; // @[Coverage map for MulAddRecFNPipe]
  wire  MulAddRecFNPipe_cov_write_addr; // @[Coverage map for MulAddRecFNPipe]
  wire  MulAddRecFNPipe_cov_write_mask; // @[Coverage map for MulAddRecFNPipe]
  wire  MulAddRecFNPipe_cov_write_en; // @[Coverage map for MulAddRecFNPipe]
  reg [29:0] MulAddRecFNPipe_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_32;
  wire  valid_stage0_shl;
  wire  valid_stage0_pad;
  wire [29:0] mulAddRecFNToRaw_preMul_sum;
  wire [29:0] mulAddRecFNToRaw_postMul_sum;
  wire [29:0] roundRawFNToRecFN_sum;
  wire  mulAddRecFNToRaw_preMul_metaAssert_wire;
  wire  mulAddRecFNToRaw_postMul_metaAssert_wire;
  wire  roundRawFNToRecFN_metaAssert_wire;
  wire  MulAddRecFNPipe_or2;
  wire  MulAddRecFNPipe_or0;
  reg  MulAddRecFNPipe_metaAssert;
  reg [31:0] _RAND_33;
  MulAddRecFNToRaw_preMul mulAddRecFNToRaw_preMul ( // @[FPU.scala 580:15]
    .io_op(mulAddRecFNToRaw_preMul_io_op),
    .io_a(mulAddRecFNToRaw_preMul_io_a),
    .io_b(mulAddRecFNToRaw_preMul_io_b),
    .io_c(mulAddRecFNToRaw_preMul_io_c),
    .io_mulAddA(mulAddRecFNToRaw_preMul_io_mulAddA),
    .io_mulAddB(mulAddRecFNToRaw_preMul_io_mulAddB),
    .io_mulAddC(mulAddRecFNToRaw_preMul_io_mulAddC),
    .io_toPostMul_isSigNaNAny(mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny),
    .io_toPostMul_isNaNAOrB(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB),
    .io_toPostMul_isInfA(mulAddRecFNToRaw_preMul_io_toPostMul_isInfA),
    .io_toPostMul_isZeroA(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA),
    .io_toPostMul_isInfB(mulAddRecFNToRaw_preMul_io_toPostMul_isInfB),
    .io_toPostMul_isZeroB(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB),
    .io_toPostMul_signProd(mulAddRecFNToRaw_preMul_io_toPostMul_signProd),
    .io_toPostMul_isNaNC(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC),
    .io_toPostMul_isInfC(mulAddRecFNToRaw_preMul_io_toPostMul_isInfC),
    .io_toPostMul_isZeroC(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC),
    .io_toPostMul_sExpSum(mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum),
    .io_toPostMul_doSubMags(mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags),
    .io_toPostMul_CIsDominant(mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant),
    .io_toPostMul_CDom_CAlignDist(mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist),
    .io_toPostMul_highAlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC),
    .io_toPostMul_bit0AlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC),
    .io_covSum(mulAddRecFNToRaw_preMul_io_covSum),
    .metaAssert(mulAddRecFNToRaw_preMul_metaAssert)
  );
  MulAddRecFNToRaw_postMul mulAddRecFNToRaw_postMul ( // @[FPU.scala 582:15]
    .io_fromPreMul_isSigNaNAny(mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny),
    .io_fromPreMul_isNaNAOrB(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB),
    .io_fromPreMul_isInfA(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA),
    .io_fromPreMul_isZeroA(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA),
    .io_fromPreMul_isInfB(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB),
    .io_fromPreMul_isZeroB(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB),
    .io_fromPreMul_signProd(mulAddRecFNToRaw_postMul_io_fromPreMul_signProd),
    .io_fromPreMul_isNaNC(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC),
    .io_fromPreMul_isInfC(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC),
    .io_fromPreMul_isZeroC(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC),
    .io_fromPreMul_sExpSum(mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum),
    .io_fromPreMul_doSubMags(mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags),
    .io_fromPreMul_CIsDominant(mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant),
    .io_fromPreMul_CDom_CAlignDist(mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist),
    .io_fromPreMul_highAlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC),
    .io_fromPreMul_bit0AlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC),
    .io_mulAddResult(mulAddRecFNToRaw_postMul_io_mulAddResult),
    .io_roundingMode(mulAddRecFNToRaw_postMul_io_roundingMode),
    .io_invalidExc(mulAddRecFNToRaw_postMul_io_invalidExc),
    .io_rawOut_isNaN(mulAddRecFNToRaw_postMul_io_rawOut_isNaN),
    .io_rawOut_isInf(mulAddRecFNToRaw_postMul_io_rawOut_isInf),
    .io_rawOut_isZero(mulAddRecFNToRaw_postMul_io_rawOut_isZero),
    .io_rawOut_sign(mulAddRecFNToRaw_postMul_io_rawOut_sign),
    .io_rawOut_sExp(mulAddRecFNToRaw_postMul_io_rawOut_sExp),
    .io_rawOut_sig(mulAddRecFNToRaw_postMul_io_rawOut_sig),
    .io_covSum(mulAddRecFNToRaw_postMul_io_covSum),
    .metaAssert(mulAddRecFNToRaw_postMul_metaAssert)
  );
  RoundRawFNToRecFN_2 roundRawFNToRecFN ( // @[FPU.scala 608:35]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_infiniteExc(roundRawFNToRecFN_io_infiniteExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundRawFNToRecFN_io_detectTininess),
    .io_out(roundRawFNToRecFN_io_out),
    .io_exceptionFlags(roundRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundRawFNToRecFN_io_covSum),
    .metaAssert(roundRawFNToRecFN_metaAssert)
  );
  assign _T_14 = mulAddRecFNToRaw_preMul_io_mulAddA * mulAddRecFNToRaw_preMul_io_mulAddB; // @[FPU.scala 590:45]
  assign mulAddResult = _T_14 + mulAddRecFNToRaw_preMul_io_mulAddC; // @[FPU.scala 591:50]
  assign io_out = roundRawFNToRecFN_io_out; // @[FPU.scala 619:23]
  assign io_exceptionFlags = roundRawFNToRecFN_io_exceptionFlags; // @[FPU.scala 620:23]
  assign mulAddRecFNToRaw_preMul_io_op = io_op; // @[FPU.scala 584:35]
  assign mulAddRecFNToRaw_preMul_io_a = io_a; // @[FPU.scala 585:35]
  assign mulAddRecFNToRaw_preMul_io_b = io_b; // @[FPU.scala 586:35]
  assign mulAddRecFNToRaw_preMul_io_c = io_c; // @[FPU.scala 587:35]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny = _T_21_isSigNaNAny; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB = _T_21_isNaNAOrB; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA = _T_21_isInfA; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA = _T_21_isZeroA; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB = _T_21_isInfB; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB = _T_21_isZeroB; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_signProd = _T_21_signProd; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC = _T_21_isNaNC; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC = _T_21_isInfC; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC = _T_21_isZeroC; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum = _T_21_sExpSum; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags = _T_21_doSubMags; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant = _T_21_CIsDominant; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist = _T_21_CDom_CAlignDist; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC = _T_21_highAlignedSigC; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC = _T_21_bit0AlignedSigC; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_mulAddResult = _T_30; // @[FPU.scala 600:46]
  assign mulAddRecFNToRaw_postMul_io_roundingMode = _T_39; // @[FPU.scala 601:46]
  assign roundRawFNToRecFN_io_invalidExc = _T_75; // @[FPU.scala 611:45]
  assign roundRawFNToRecFN_io_infiniteExc = 1'h0; // @[FPU.scala 617:38]
  assign roundRawFNToRecFN_io_in_isNaN = _T_84_isNaN; // @[FPU.scala 612:45]
  assign roundRawFNToRecFN_io_in_isInf = _T_84_isInf; // @[FPU.scala 612:45]
  assign roundRawFNToRecFN_io_in_isZero = _T_84_isZero; // @[FPU.scala 612:45]
  assign roundRawFNToRecFN_io_in_sign = _T_84_sign; // @[FPU.scala 612:45]
  assign roundRawFNToRecFN_io_in_sExp = _T_84_sExp; // @[FPU.scala 612:45]
  assign roundRawFNToRecFN_io_in_sig = _T_84_sig; // @[FPU.scala 612:45]
  assign roundRawFNToRecFN_io_roundingMode = _T_93; // @[FPU.scala 613:45]
  assign roundRawFNToRecFN_io_detectTininess = _T_102; // @[FPU.scala 614:45]
  assign MulAddRecFNPipe_cov_read_addr = MulAddRecFNPipe_state;
  assign MulAddRecFNPipe_cov_read_data = MulAddRecFNPipe_cov[MulAddRecFNPipe_cov_read_addr]; // @[Coverage map for MulAddRecFNPipe]
  assign MulAddRecFNPipe_cov_write_data = 1'h1;
  assign MulAddRecFNPipe_cov_write_addr = MulAddRecFNPipe_state;
  assign MulAddRecFNPipe_cov_write_mask = 1'h1;
  assign MulAddRecFNPipe_cov_write_en = 1'h1;
  assign valid_stage0_shl = valid_stage0;
  assign valid_stage0_pad = valid_stage0_shl;
  assign mulAddRecFNToRaw_preMul_sum = MulAddRecFNPipe_covSum + mulAddRecFNToRaw_preMul_io_covSum;
  assign mulAddRecFNToRaw_postMul_sum = mulAddRecFNToRaw_preMul_sum + mulAddRecFNToRaw_postMul_io_covSum;
  assign roundRawFNToRecFN_sum = mulAddRecFNToRaw_postMul_sum + roundRawFNToRecFN_io_covSum;
  assign io_covSum = roundRawFNToRecFN_sum;
  assign mulAddRecFNToRaw_preMul_metaAssert_wire = mulAddRecFNToRaw_preMul_metaAssert;
  assign mulAddRecFNToRaw_postMul_metaAssert_wire = mulAddRecFNToRaw_postMul_metaAssert;
  assign roundRawFNToRecFN_metaAssert_wire = roundRawFNToRecFN_metaAssert;
  assign MulAddRecFNPipe_or2 = mulAddRecFNToRaw_postMul_metaAssert_wire | roundRawFNToRecFN_metaAssert_wire;
  assign MulAddRecFNPipe_or0 = mulAddRecFNToRaw_preMul_metaAssert_wire | MulAddRecFNPipe_or2;
  assign metaAssert = MulAddRecFNPipe_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_21_isSigNaNAny = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_21_isNaNAOrB = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_21_isInfA = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_21_isZeroA = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_21_isInfB = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_21_isZeroB = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_21_signProd = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_21_isNaNC = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_21_isInfC = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_21_isZeroC = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_21_sExpSum = _RAND_10[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_21_doSubMags = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_21_CIsDominant = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_21_CDom_CAlignDist = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_21_highAlignedSigC = _RAND_14[25:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_21_bit0AlignedSigC = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {2{`RANDOM}};
  _T_30 = _RAND_16[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_39 = _RAND_17[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  roundingMode_stage0 = _RAND_18[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  detectTininess_stage0 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  valid_stage0 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_75 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_84_isNaN = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_84_isInf = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_84_isZero = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_84_sign = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_84_sExp = _RAND_26[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_84_sig = _RAND_27[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_93 = _RAND_28[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_102 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  MulAddRecFNPipe_state = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    MulAddRecFNPipe_cov[initvar] = _RAND_31[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  MulAddRecFNPipe_covSum = _RAND_32[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  MulAddRecFNPipe_metaAssert = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      _T_21_isSigNaNAny <= 1'h0;
    end else if (io_validin) begin
      _T_21_isSigNaNAny <= mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny;
    end
    if (metaReset) begin
      _T_21_isNaNAOrB <= 1'h0;
    end else if (io_validin) begin
      _T_21_isNaNAOrB <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB;
    end
    if (metaReset) begin
      _T_21_isInfA <= 1'h0;
    end else if (io_validin) begin
      _T_21_isInfA <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfA;
    end
    if (metaReset) begin
      _T_21_isZeroA <= 1'h0;
    end else if (io_validin) begin
      _T_21_isZeroA <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA;
    end
    if (metaReset) begin
      _T_21_isInfB <= 1'h0;
    end else if (io_validin) begin
      _T_21_isInfB <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfB;
    end
    if (metaReset) begin
      _T_21_isZeroB <= 1'h0;
    end else if (io_validin) begin
      _T_21_isZeroB <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB;
    end
    if (metaReset) begin
      _T_21_signProd <= 1'h0;
    end else if (io_validin) begin
      _T_21_signProd <= mulAddRecFNToRaw_preMul_io_toPostMul_signProd;
    end
    if (metaReset) begin
      _T_21_isNaNC <= 1'h0;
    end else if (io_validin) begin
      _T_21_isNaNC <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC;
    end
    if (metaReset) begin
      _T_21_isInfC <= 1'h0;
    end else if (io_validin) begin
      _T_21_isInfC <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfC;
    end
    if (metaReset) begin
      _T_21_isZeroC <= 1'h0;
    end else if (io_validin) begin
      _T_21_isZeroC <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC;
    end
    if (metaReset) begin
      _T_21_sExpSum <= 10'h0;
    end else if (io_validin) begin
      _T_21_sExpSum <= mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum;
    end
    if (metaReset) begin
      _T_21_doSubMags <= 1'h0;
    end else if (io_validin) begin
      _T_21_doSubMags <= mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags;
    end
    if (metaReset) begin
      _T_21_CIsDominant <= 1'h0;
    end else if (io_validin) begin
      _T_21_CIsDominant <= mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant;
    end
    if (metaReset) begin
      _T_21_CDom_CAlignDist <= 5'h0;
    end else if (io_validin) begin
      _T_21_CDom_CAlignDist <= mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist;
    end
    if (metaReset) begin
      _T_21_highAlignedSigC <= 26'h0;
    end else if (io_validin) begin
      _T_21_highAlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC;
    end
    if (metaReset) begin
      _T_21_bit0AlignedSigC <= 1'h0;
    end else if (io_validin) begin
      _T_21_bit0AlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC;
    end
    if (metaReset) begin
      _T_30 <= 49'h0;
    end else if (io_validin) begin
      _T_30 <= mulAddResult;
    end
    if (metaReset) begin
      _T_39 <= 3'h0;
    end else if (io_validin) begin
      _T_39 <= io_roundingMode;
    end
    if (metaReset) begin
      roundingMode_stage0 <= 3'h0;
    end else if (io_validin) begin
      roundingMode_stage0 <= io_roundingMode;
    end
    if (metaReset) begin
      detectTininess_stage0 <= 1'h0;
    end else begin
      detectTininess_stage0 <= io_validin | detectTininess_stage0;
    end
    if (metaReset) begin
      valid_stage0 <= 1'h0;
    end else if (reset) begin
      valid_stage0 <= 1'h0;
    end else begin
      valid_stage0 <= io_validin;
    end
    if (metaReset) begin
      _T_75 <= 1'h0;
    end else if (valid_stage0) begin
      _T_75 <= mulAddRecFNToRaw_postMul_io_invalidExc;
    end
    if (metaReset) begin
      _T_84_isNaN <= 1'h0;
    end else if (valid_stage0) begin
      _T_84_isNaN <= mulAddRecFNToRaw_postMul_io_rawOut_isNaN;
    end
    if (metaReset) begin
      _T_84_isInf <= 1'h0;
    end else if (valid_stage0) begin
      _T_84_isInf <= mulAddRecFNToRaw_postMul_io_rawOut_isInf;
    end
    if (metaReset) begin
      _T_84_isZero <= 1'h0;
    end else if (valid_stage0) begin
      _T_84_isZero <= mulAddRecFNToRaw_postMul_io_rawOut_isZero;
    end
    if (metaReset) begin
      _T_84_sign <= 1'h0;
    end else if (valid_stage0) begin
      _T_84_sign <= mulAddRecFNToRaw_postMul_io_rawOut_sign;
    end
    if (metaReset) begin
      _T_84_sExp <= 10'h0;
    end else if (valid_stage0) begin
      _T_84_sExp <= mulAddRecFNToRaw_postMul_io_rawOut_sExp;
    end
    if (metaReset) begin
      _T_84_sig <= 27'h0;
    end else if (valid_stage0) begin
      _T_84_sig <= mulAddRecFNToRaw_postMul_io_rawOut_sig;
    end
    if (metaReset) begin
      _T_93 <= 3'h0;
    end else if (valid_stage0) begin
      _T_93 <= roundingMode_stage0;
    end
    if (metaReset) begin
      _T_102 <= 1'h0;
    end else if (valid_stage0) begin
      _T_102 <= detectTininess_stage0;
    end
    MulAddRecFNPipe_state <= valid_stage0_pad;
    if (!(MulAddRecFNPipe_cov_read_data)) begin
      MulAddRecFNPipe_covSum <= MulAddRecFNPipe_covSum + 1'h1;
    end
    if (metaReset) begin
      MulAddRecFNPipe_metaAssert <= 1'h0;
    end else begin
      MulAddRecFNPipe_metaAssert <= MulAddRecFNPipe_metaAssert | MulAddRecFNPipe_or0;
    end
  end
  always @(posedge clock) begin
    if(MulAddRecFNPipe_cov_write_en & MulAddRecFNPipe_cov_write_mask) begin
      MulAddRecFNPipe_cov[MulAddRecFNPipe_cov_write_addr] <= MulAddRecFNPipe_cov_write_data; // @[Coverage map for MulAddRecFNPipe]
    end
  end
endmodule
module CompareRecFN(
  input  [64:0] io_a,
  input  [64:0] io_b,
  input         io_signaling,
  output        io_lt,
  output        io_eq,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  rawA_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_15; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawA_isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawA_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawA_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] rawA_sig; // @[Cat.scala 30:58]
  wire  rawB_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_32; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawB_isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawB_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawB_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] rawB_sig; // @[Cat.scala 30:58]
  wire  ordered; // @[CompareRecFN.scala 57:32]
  wire  bothInfs; // @[CompareRecFN.scala 58:33]
  wire  bothZeros; // @[CompareRecFN.scala 59:33]
  wire  eqExps; // @[CompareRecFN.scala 60:29]
  wire  _T_47; // @[CompareRecFN.scala 62:20]
  wire  _T_48; // @[CompareRecFN.scala 62:57]
  wire  _T_49; // @[CompareRecFN.scala 62:44]
  wire  common_ltMags; // @[CompareRecFN.scala 62:33]
  wire  _T_50; // @[CompareRecFN.scala 63:45]
  wire  common_eqMags; // @[CompareRecFN.scala 63:32]
  wire  _T_53; // @[CompareRecFN.scala 67:25]
  wire  _T_56; // @[CompareRecFN.scala 69:35]
  wire  _T_58; // @[CompareRecFN.scala 69:54]
  wire  _T_60; // @[CompareRecFN.scala 70:41]
  wire  _T_61; // @[CompareRecFN.scala 69:74]
  wire  _T_62; // @[CompareRecFN.scala 68:30]
  wire  _T_63; // @[CompareRecFN.scala 67:41]
  wire  ordered_lt; // @[CompareRecFN.scala 66:21]
  wire  _T_64; // @[CompareRecFN.scala 72:34]
  wire  _T_65; // @[CompareRecFN.scala 72:62]
  wire  _T_66; // @[CompareRecFN.scala 72:49]
  wire  ordered_eq; // @[CompareRecFN.scala 72:19]
  wire  _T_69; // @[common.scala 81:46]
  wire  _T_72; // @[common.scala 81:46]
  wire  _T_73; // @[CompareRecFN.scala 75:32]
  wire  _T_75; // @[CompareRecFN.scala 76:27]
  wire  invalid; // @[CompareRecFN.scala 75:58]
  wire [29:0] CompareRecFN_covSum;
  assign rawA_isZero = io_a[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_15 = io_a[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawA_isNaN = _T_15 & io_a[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawA_isInf = _T_15 & ~io_a[61]; // @[rawFloatFromRecFN.scala 56:33]
  assign rawA_sign = io_a[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawA_sExp = {1'b0,$signed(io_a[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawA_sig = {1'h0,~rawA_isZero,io_a[51:0]}; // @[Cat.scala 30:58]
  assign rawB_isZero = io_b[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_32 = io_b[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawB_isNaN = _T_32 & io_b[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawB_isInf = _T_32 & ~io_b[61]; // @[rawFloatFromRecFN.scala 56:33]
  assign rawB_sign = io_b[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawB_sExp = {1'b0,$signed(io_b[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawB_sig = {1'h0,~rawB_isZero,io_b[51:0]}; // @[Cat.scala 30:58]
  assign ordered = ~rawA_isNaN & ~rawB_isNaN; // @[CompareRecFN.scala 57:32]
  assign bothInfs = rawA_isInf & rawB_isInf; // @[CompareRecFN.scala 58:33]
  assign bothZeros = rawA_isZero & rawB_isZero; // @[CompareRecFN.scala 59:33]
  assign eqExps = $signed(rawA_sExp) == $signed(rawB_sExp); // @[CompareRecFN.scala 60:29]
  assign _T_47 = $signed(rawA_sExp) < $signed(rawB_sExp); // @[CompareRecFN.scala 62:20]
  assign _T_48 = rawA_sig < rawB_sig; // @[CompareRecFN.scala 62:57]
  assign _T_49 = eqExps & _T_48; // @[CompareRecFN.scala 62:44]
  assign common_ltMags = _T_47 | _T_49; // @[CompareRecFN.scala 62:33]
  assign _T_50 = rawA_sig == rawB_sig; // @[CompareRecFN.scala 63:45]
  assign common_eqMags = eqExps & _T_50; // @[CompareRecFN.scala 63:32]
  assign _T_53 = rawA_sign & ~rawB_sign; // @[CompareRecFN.scala 67:25]
  assign _T_56 = rawA_sign & ~common_ltMags; // @[CompareRecFN.scala 69:35]
  assign _T_58 = _T_56 & ~common_eqMags; // @[CompareRecFN.scala 69:54]
  assign _T_60 = ~rawB_sign & common_ltMags; // @[CompareRecFN.scala 70:41]
  assign _T_61 = _T_58 | _T_60; // @[CompareRecFN.scala 69:74]
  assign _T_62 = ~bothInfs & _T_61; // @[CompareRecFN.scala 68:30]
  assign _T_63 = _T_53 | _T_62; // @[CompareRecFN.scala 67:41]
  assign ordered_lt = ~bothZeros & _T_63; // @[CompareRecFN.scala 66:21]
  assign _T_64 = rawA_sign == rawB_sign; // @[CompareRecFN.scala 72:34]
  assign _T_65 = bothInfs | common_eqMags; // @[CompareRecFN.scala 72:62]
  assign _T_66 = _T_64 & _T_65; // @[CompareRecFN.scala 72:49]
  assign ordered_eq = bothZeros | _T_66; // @[CompareRecFN.scala 72:19]
  assign _T_69 = rawA_isNaN & ~rawA_sig[51]; // @[common.scala 81:46]
  assign _T_72 = rawB_isNaN & ~rawB_sig[51]; // @[common.scala 81:46]
  assign _T_73 = _T_69 | _T_72; // @[CompareRecFN.scala 75:32]
  assign _T_75 = io_signaling & ~ordered; // @[CompareRecFN.scala 76:27]
  assign invalid = _T_73 | _T_75; // @[CompareRecFN.scala 75:58]
  assign io_lt = ordered & ordered_lt; // @[CompareRecFN.scala 78:11]
  assign io_eq = ordered & ordered_eq; // @[CompareRecFN.scala 79:11]
  assign io_exceptionFlags = {invalid,4'h0}; // @[CompareRecFN.scala 81:23]
  assign CompareRecFN_covSum = 30'h0;
  assign io_covSum = CompareRecFN_covSum;
  assign metaAssert = 1'h0;
endmodule
module RecFNToIN(
  input  [64:0] io_in,
  input  [2:0]  io_roundingMode,
  input         io_signedOut,
  output [63:0] io_out,
  output [2:0]  io_intExceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  rawIn_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_13; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawIn_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawIn_isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawIn_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawIn_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] rawIn_sig; // @[Cat.scala 30:58]
  wire  magGeOne; // @[RecFNToIN.scala 58:30]
  wire [10:0] posExp; // @[RecFNToIN.scala 59:28]
  wire  _T_28; // @[RecFNToIN.scala 60:48]
  wire  magJustBelowOne; // @[RecFNToIN.scala 60:38]
  wire  roundingMode_near_even; // @[RecFNToIN.scala 64:53]
  wire  roundingMode_min; // @[RecFNToIN.scala 67:53]
  wire  roundingMode_max; // @[RecFNToIN.scala 68:53]
  wire  roundingMode_near_maxMag; // @[RecFNToIN.scala 69:53]
  wire [52:0] _T_32; // @[Cat.scala 30:58]
  wire [5:0] _T_34; // @[RecFNToIN.scala 81:16]
  wire [115:0] _GEN_0; // @[RecFNToIN.scala 80:50]
  wire [115:0] shiftedSig; // @[RecFNToIN.scala 80:50]
  wire  _T_37; // @[RecFNToIN.scala 86:69]
  wire [65:0] alignedSig; // @[Cat.scala 30:58]
  wire [63:0] unroundedInt; // @[RecFNToIN.scala 87:54]
  wire  _T_40; // @[RecFNToIN.scala 89:57]
  wire  common_inexact; // @[RecFNToIN.scala 89:29]
  wire  _T_44; // @[RecFNToIN.scala 91:46]
  wire  _T_47; // @[RecFNToIN.scala 91:71]
  wire  _T_48; // @[RecFNToIN.scala 91:51]
  wire  _T_49; // @[RecFNToIN.scala 91:25]
  wire  _T_52; // @[RecFNToIN.scala 92:26]
  wire  roundIncr_near_even; // @[RecFNToIN.scala 91:78]
  wire  _T_54; // @[RecFNToIN.scala 93:43]
  wire  roundIncr_near_maxMag; // @[RecFNToIN.scala 93:61]
  wire  _T_55; // @[RecFNToIN.scala 95:35]
  wire  _T_56; // @[RecFNToIN.scala 96:35]
  wire  _T_57; // @[RecFNToIN.scala 95:72]
  wire  _T_58; // @[RecFNToIN.scala 97:52]
  wire  _T_59; // @[RecFNToIN.scala 97:35]
  wire  _T_60; // @[RecFNToIN.scala 96:72]
  wire  _T_62; // @[RecFNToIN.scala 98:52]
  wire  _T_63; // @[RecFNToIN.scala 98:35]
  wire  roundIncr; // @[RecFNToIN.scala 97:72]
  wire [63:0] complUnroundedInt; // @[RecFNToIN.scala 99:32]
  wire  _T_65; // @[RecFNToIN.scala 101:23]
  wire [63:0] _T_67; // @[RecFNToIN.scala 102:31]
  wire [63:0] roundedInt; // @[RecFNToIN.scala 101:12]
  wire  magGeOne_atOverflowEdge; // @[RecFNToIN.scala 106:43]
  wire  _T_70; // @[RecFNToIN.scala 109:56]
  wire  roundCarryBut2; // @[RecFNToIN.scala 109:61]
  wire  _T_71; // @[RecFNToIN.scala 112:21]
  wire  _T_73; // @[RecFNToIN.scala 116:60]
  wire  _T_74; // @[RecFNToIN.scala 116:64]
  wire  _T_75; // @[RecFNToIN.scala 115:49]
  wire  _T_76; // @[RecFNToIN.scala 118:38]
  wire  _T_77; // @[RecFNToIN.scala 118:62]
  wire  _T_78; // @[RecFNToIN.scala 117:49]
  wire  _T_79; // @[RecFNToIN.scala 114:24]
  wire  _T_81; // @[RecFNToIN.scala 121:50]
  wire  _T_82; // @[RecFNToIN.scala 122:57]
  wire  _T_83; // @[RecFNToIN.scala 120:32]
  wire  _T_84; // @[RecFNToIN.scala 113:20]
  wire  _T_85; // @[RecFNToIN.scala 112:40]
  wire  _T_87; // @[RecFNToIN.scala 124:28]
  wire  _T_88; // @[RecFNToIN.scala 124:42]
  wire  common_overflow; // @[RecFNToIN.scala 111:12]
  wire  invalidExc; // @[RecFNToIN.scala 129:34]
  wire  overflow; // @[RecFNToIN.scala 130:33]
  wire  _T_92; // @[RecFNToIN.scala 131:33]
  wire  inexact; // @[RecFNToIN.scala 131:54]
  wire  excSign; // @[RecFNToIN.scala 133:33]
  wire  _T_94; // @[RecFNToIN.scala 135:27]
  wire [63:0] _T_95; // @[RecFNToIN.scala 135:12]
  wire [62:0] _T_97; // @[RecFNToIN.scala 139:12]
  wire [63:0] _GEN_1; // @[RecFNToIN.scala 138:11]
  wire [63:0] excOut; // @[RecFNToIN.scala 138:11]
  wire  _T_98; // @[RecFNToIN.scala 141:30]
  wire [1:0] _T_100; // @[Cat.scala 30:58]
  wire [29:0] RecFNToIN_covSum;
  assign rawIn_isZero = io_in[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_13 = io_in[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawIn_isNaN = _T_13 & io_in[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawIn_isInf = _T_13 & ~io_in[61]; // @[rawFloatFromRecFN.scala 56:33]
  assign rawIn_sign = io_in[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawIn_sExp = {1'b0,$signed(io_in[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawIn_sig = {1'h0,~rawIn_isZero,io_in[51:0]}; // @[Cat.scala 30:58]
  assign magGeOne = rawIn_sExp[11]; // @[RecFNToIN.scala 58:30]
  assign posExp = rawIn_sExp[10:0]; // @[RecFNToIN.scala 59:28]
  assign _T_28 = ~posExp == 11'h0; // @[RecFNToIN.scala 60:48]
  assign magJustBelowOne = ~magGeOne & _T_28; // @[RecFNToIN.scala 60:38]
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RecFNToIN.scala 64:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RecFNToIN.scala 67:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RecFNToIN.scala 68:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RecFNToIN.scala 69:53]
  assign _T_32 = {magGeOne,rawIn_sig[51:0]}; // @[Cat.scala 30:58]
  assign _T_34 = magGeOne ? rawIn_sExp[5:0] : 6'h0; // @[RecFNToIN.scala 81:16]
  assign _GEN_0 = {{63'd0}, _T_32}; // @[RecFNToIN.scala 80:50]
  assign shiftedSig = _GEN_0 << _T_34; // @[RecFNToIN.scala 80:50]
  assign _T_37 = shiftedSig[50:0] != 51'h0; // @[RecFNToIN.scala 86:69]
  assign alignedSig = {shiftedSig[115:51],_T_37}; // @[Cat.scala 30:58]
  assign unroundedInt = alignedSig[65:2]; // @[RecFNToIN.scala 87:54]
  assign _T_40 = alignedSig[1:0] != 2'h0; // @[RecFNToIN.scala 89:57]
  assign common_inexact = magGeOne ? _T_40 : ~rawIn_isZero; // @[RecFNToIN.scala 89:29]
  assign _T_44 = ~alignedSig[2:1] == 2'h0; // @[RecFNToIN.scala 91:46]
  assign _T_47 = ~alignedSig[1:0] == 2'h0; // @[RecFNToIN.scala 91:71]
  assign _T_48 = _T_44 | _T_47; // @[RecFNToIN.scala 91:51]
  assign _T_49 = magGeOne & _T_48; // @[RecFNToIN.scala 91:25]
  assign _T_52 = magJustBelowOne & _T_40; // @[RecFNToIN.scala 92:26]
  assign roundIncr_near_even = _T_49 | _T_52; // @[RecFNToIN.scala 91:78]
  assign _T_54 = magGeOne & alignedSig[1]; // @[RecFNToIN.scala 93:43]
  assign roundIncr_near_maxMag = _T_54 | magJustBelowOne; // @[RecFNToIN.scala 93:61]
  assign _T_55 = roundingMode_near_even & roundIncr_near_even; // @[RecFNToIN.scala 95:35]
  assign _T_56 = roundingMode_near_maxMag & roundIncr_near_maxMag; // @[RecFNToIN.scala 96:35]
  assign _T_57 = _T_55 | _T_56; // @[RecFNToIN.scala 95:72]
  assign _T_58 = rawIn_sign & common_inexact; // @[RecFNToIN.scala 97:52]
  assign _T_59 = roundingMode_min & _T_58; // @[RecFNToIN.scala 97:35]
  assign _T_60 = _T_57 | _T_59; // @[RecFNToIN.scala 96:72]
  assign _T_62 = ~rawIn_sign & common_inexact; // @[RecFNToIN.scala 98:52]
  assign _T_63 = roundingMode_max & _T_62; // @[RecFNToIN.scala 98:35]
  assign roundIncr = _T_60 | _T_63; // @[RecFNToIN.scala 97:72]
  assign complUnroundedInt = rawIn_sign ? ~unroundedInt : unroundedInt; // @[RecFNToIN.scala 99:32]
  assign _T_65 = roundIncr ^ rawIn_sign; // @[RecFNToIN.scala 101:23]
  assign _T_67 = complUnroundedInt + 64'h1; // @[RecFNToIN.scala 102:31]
  assign roundedInt = _T_65 ? _T_67 : complUnroundedInt; // @[RecFNToIN.scala 101:12]
  assign magGeOne_atOverflowEdge = posExp == 11'h3f; // @[RecFNToIN.scala 106:43]
  assign _T_70 = ~unroundedInt[61:0] == 62'h0; // @[RecFNToIN.scala 109:56]
  assign roundCarryBut2 = _T_70 & roundIncr; // @[RecFNToIN.scala 109:61]
  assign _T_71 = posExp >= 11'h40; // @[RecFNToIN.scala 112:21]
  assign _T_73 = unroundedInt[62:0] != 63'h0; // @[RecFNToIN.scala 116:60]
  assign _T_74 = _T_73 | roundIncr; // @[RecFNToIN.scala 116:64]
  assign _T_75 = magGeOne_atOverflowEdge & _T_74; // @[RecFNToIN.scala 115:49]
  assign _T_76 = posExp == 11'h3e; // @[RecFNToIN.scala 118:38]
  assign _T_77 = _T_76 & roundCarryBut2; // @[RecFNToIN.scala 118:62]
  assign _T_78 = magGeOne_atOverflowEdge | _T_77; // @[RecFNToIN.scala 117:49]
  assign _T_79 = rawIn_sign ? _T_75 : _T_78; // @[RecFNToIN.scala 114:24]
  assign _T_81 = magGeOne_atOverflowEdge & unroundedInt[62]; // @[RecFNToIN.scala 121:50]
  assign _T_82 = _T_81 & roundCarryBut2; // @[RecFNToIN.scala 122:57]
  assign _T_83 = rawIn_sign | _T_82; // @[RecFNToIN.scala 120:32]
  assign _T_84 = io_signedOut ? _T_79 : _T_83; // @[RecFNToIN.scala 113:20]
  assign _T_85 = _T_71 | _T_84; // @[RecFNToIN.scala 112:40]
  assign _T_87 = ~io_signedOut & rawIn_sign; // @[RecFNToIN.scala 124:28]
  assign _T_88 = _T_87 & roundIncr; // @[RecFNToIN.scala 124:42]
  assign common_overflow = magGeOne ? _T_85 : _T_88; // @[RecFNToIN.scala 111:12]
  assign invalidExc = rawIn_isNaN | rawIn_isInf; // @[RecFNToIN.scala 129:34]
  assign overflow = ~invalidExc & common_overflow; // @[RecFNToIN.scala 130:33]
  assign _T_92 = ~invalidExc & ~common_overflow; // @[RecFNToIN.scala 131:33]
  assign inexact = _T_92 & common_inexact; // @[RecFNToIN.scala 131:54]
  assign excSign = ~rawIn_isNaN & rawIn_sign; // @[RecFNToIN.scala 133:33]
  assign _T_94 = io_signedOut == excSign; // @[RecFNToIN.scala 135:27]
  assign _T_95 = _T_94 ? 64'h8000000000000000 : 64'h0; // @[RecFNToIN.scala 135:12]
  assign _T_97 = excSign ? 63'h0 : 63'h7fffffffffffffff; // @[RecFNToIN.scala 139:12]
  assign _GEN_1 = {{1'd0}, _T_97}; // @[RecFNToIN.scala 138:11]
  assign excOut = _T_95 | _GEN_1; // @[RecFNToIN.scala 138:11]
  assign _T_98 = invalidExc | common_overflow; // @[RecFNToIN.scala 141:30]
  assign _T_100 = {invalidExc,overflow}; // @[Cat.scala 30:58]
  assign io_out = _T_98 ? excOut : roundedInt; // @[RecFNToIN.scala 141:12]
  assign io_intExceptionFlags = {_T_100,inexact}; // @[RecFNToIN.scala 142:26]
  assign RecFNToIN_covSum = 30'h0;
  assign io_covSum = RecFNToIN_covSum;
  assign metaAssert = 1'h0;
endmodule
module RecFNToIN_1(
  input  [64:0] io_in,
  input  [2:0]  io_roundingMode,
  input         io_signedOut,
  output [2:0]  io_intExceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  rawIn_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_13; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawIn_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawIn_isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawIn_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawIn_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] rawIn_sig; // @[Cat.scala 30:58]
  wire  magGeOne; // @[RecFNToIN.scala 58:30]
  wire [10:0] posExp; // @[RecFNToIN.scala 59:28]
  wire  _T_28; // @[RecFNToIN.scala 60:48]
  wire  magJustBelowOne; // @[RecFNToIN.scala 60:38]
  wire  roundingMode_near_even; // @[RecFNToIN.scala 64:53]
  wire  roundingMode_min; // @[RecFNToIN.scala 67:53]
  wire  roundingMode_max; // @[RecFNToIN.scala 68:53]
  wire  roundingMode_near_maxMag; // @[RecFNToIN.scala 69:53]
  wire [52:0] _T_32; // @[Cat.scala 30:58]
  wire [4:0] _T_34; // @[RecFNToIN.scala 81:16]
  wire [83:0] _GEN_0; // @[RecFNToIN.scala 80:50]
  wire [83:0] shiftedSig; // @[RecFNToIN.scala 80:50]
  wire  _T_37; // @[RecFNToIN.scala 86:69]
  wire [33:0] alignedSig; // @[Cat.scala 30:58]
  wire [31:0] unroundedInt; // @[RecFNToIN.scala 87:54]
  wire  _T_40; // @[RecFNToIN.scala 89:57]
  wire  common_inexact; // @[RecFNToIN.scala 89:29]
  wire  _T_44; // @[RecFNToIN.scala 91:46]
  wire  _T_47; // @[RecFNToIN.scala 91:71]
  wire  _T_48; // @[RecFNToIN.scala 91:51]
  wire  _T_49; // @[RecFNToIN.scala 91:25]
  wire  _T_52; // @[RecFNToIN.scala 92:26]
  wire  roundIncr_near_even; // @[RecFNToIN.scala 91:78]
  wire  _T_54; // @[RecFNToIN.scala 93:43]
  wire  roundIncr_near_maxMag; // @[RecFNToIN.scala 93:61]
  wire  _T_55; // @[RecFNToIN.scala 95:35]
  wire  _T_56; // @[RecFNToIN.scala 96:35]
  wire  _T_57; // @[RecFNToIN.scala 95:72]
  wire  _T_58; // @[RecFNToIN.scala 97:52]
  wire  _T_59; // @[RecFNToIN.scala 97:35]
  wire  _T_60; // @[RecFNToIN.scala 96:72]
  wire  _T_62; // @[RecFNToIN.scala 98:52]
  wire  _T_63; // @[RecFNToIN.scala 98:35]
  wire  roundIncr; // @[RecFNToIN.scala 97:72]
  wire  magGeOne_atOverflowEdge; // @[RecFNToIN.scala 106:43]
  wire  _T_70; // @[RecFNToIN.scala 109:56]
  wire  roundCarryBut2; // @[RecFNToIN.scala 109:61]
  wire  _T_71; // @[RecFNToIN.scala 112:21]
  wire  _T_73; // @[RecFNToIN.scala 116:60]
  wire  _T_74; // @[RecFNToIN.scala 116:64]
  wire  _T_75; // @[RecFNToIN.scala 115:49]
  wire  _T_76; // @[RecFNToIN.scala 118:38]
  wire  _T_77; // @[RecFNToIN.scala 118:62]
  wire  _T_78; // @[RecFNToIN.scala 117:49]
  wire  _T_79; // @[RecFNToIN.scala 114:24]
  wire  _T_81; // @[RecFNToIN.scala 121:50]
  wire  _T_82; // @[RecFNToIN.scala 122:57]
  wire  _T_83; // @[RecFNToIN.scala 120:32]
  wire  _T_84; // @[RecFNToIN.scala 113:20]
  wire  _T_85; // @[RecFNToIN.scala 112:40]
  wire  _T_87; // @[RecFNToIN.scala 124:28]
  wire  _T_88; // @[RecFNToIN.scala 124:42]
  wire  common_overflow; // @[RecFNToIN.scala 111:12]
  wire  invalidExc; // @[RecFNToIN.scala 129:34]
  wire  overflow; // @[RecFNToIN.scala 130:33]
  wire  _T_92; // @[RecFNToIN.scala 131:33]
  wire  inexact; // @[RecFNToIN.scala 131:54]
  wire [1:0] _T_100; // @[Cat.scala 30:58]
  wire [29:0] RecFNToIN_1_covSum;
  assign rawIn_isZero = io_in[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_13 = io_in[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawIn_isNaN = _T_13 & io_in[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawIn_isInf = _T_13 & ~io_in[61]; // @[rawFloatFromRecFN.scala 56:33]
  assign rawIn_sign = io_in[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawIn_sExp = {1'b0,$signed(io_in[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawIn_sig = {1'h0,~rawIn_isZero,io_in[51:0]}; // @[Cat.scala 30:58]
  assign magGeOne = rawIn_sExp[11]; // @[RecFNToIN.scala 58:30]
  assign posExp = rawIn_sExp[10:0]; // @[RecFNToIN.scala 59:28]
  assign _T_28 = ~posExp == 11'h0; // @[RecFNToIN.scala 60:48]
  assign magJustBelowOne = ~magGeOne & _T_28; // @[RecFNToIN.scala 60:38]
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RecFNToIN.scala 64:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RecFNToIN.scala 67:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RecFNToIN.scala 68:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RecFNToIN.scala 69:53]
  assign _T_32 = {magGeOne,rawIn_sig[51:0]}; // @[Cat.scala 30:58]
  assign _T_34 = magGeOne ? rawIn_sExp[4:0] : 5'h0; // @[RecFNToIN.scala 81:16]
  assign _GEN_0 = {{31'd0}, _T_32}; // @[RecFNToIN.scala 80:50]
  assign shiftedSig = _GEN_0 << _T_34; // @[RecFNToIN.scala 80:50]
  assign _T_37 = shiftedSig[50:0] != 51'h0; // @[RecFNToIN.scala 86:69]
  assign alignedSig = {shiftedSig[83:51],_T_37}; // @[Cat.scala 30:58]
  assign unroundedInt = alignedSig[33:2]; // @[RecFNToIN.scala 87:54]
  assign _T_40 = alignedSig[1:0] != 2'h0; // @[RecFNToIN.scala 89:57]
  assign common_inexact = magGeOne ? _T_40 : ~rawIn_isZero; // @[RecFNToIN.scala 89:29]
  assign _T_44 = ~alignedSig[2:1] == 2'h0; // @[RecFNToIN.scala 91:46]
  assign _T_47 = ~alignedSig[1:0] == 2'h0; // @[RecFNToIN.scala 91:71]
  assign _T_48 = _T_44 | _T_47; // @[RecFNToIN.scala 91:51]
  assign _T_49 = magGeOne & _T_48; // @[RecFNToIN.scala 91:25]
  assign _T_52 = magJustBelowOne & _T_40; // @[RecFNToIN.scala 92:26]
  assign roundIncr_near_even = _T_49 | _T_52; // @[RecFNToIN.scala 91:78]
  assign _T_54 = magGeOne & alignedSig[1]; // @[RecFNToIN.scala 93:43]
  assign roundIncr_near_maxMag = _T_54 | magJustBelowOne; // @[RecFNToIN.scala 93:61]
  assign _T_55 = roundingMode_near_even & roundIncr_near_even; // @[RecFNToIN.scala 95:35]
  assign _T_56 = roundingMode_near_maxMag & roundIncr_near_maxMag; // @[RecFNToIN.scala 96:35]
  assign _T_57 = _T_55 | _T_56; // @[RecFNToIN.scala 95:72]
  assign _T_58 = rawIn_sign & common_inexact; // @[RecFNToIN.scala 97:52]
  assign _T_59 = roundingMode_min & _T_58; // @[RecFNToIN.scala 97:35]
  assign _T_60 = _T_57 | _T_59; // @[RecFNToIN.scala 96:72]
  assign _T_62 = ~rawIn_sign & common_inexact; // @[RecFNToIN.scala 98:52]
  assign _T_63 = roundingMode_max & _T_62; // @[RecFNToIN.scala 98:35]
  assign roundIncr = _T_60 | _T_63; // @[RecFNToIN.scala 97:72]
  assign magGeOne_atOverflowEdge = posExp == 11'h1f; // @[RecFNToIN.scala 106:43]
  assign _T_70 = ~unroundedInt[29:0] == 30'h0; // @[RecFNToIN.scala 109:56]
  assign roundCarryBut2 = _T_70 & roundIncr; // @[RecFNToIN.scala 109:61]
  assign _T_71 = posExp >= 11'h20; // @[RecFNToIN.scala 112:21]
  assign _T_73 = unroundedInt[30:0] != 31'h0; // @[RecFNToIN.scala 116:60]
  assign _T_74 = _T_73 | roundIncr; // @[RecFNToIN.scala 116:64]
  assign _T_75 = magGeOne_atOverflowEdge & _T_74; // @[RecFNToIN.scala 115:49]
  assign _T_76 = posExp == 11'h1e; // @[RecFNToIN.scala 118:38]
  assign _T_77 = _T_76 & roundCarryBut2; // @[RecFNToIN.scala 118:62]
  assign _T_78 = magGeOne_atOverflowEdge | _T_77; // @[RecFNToIN.scala 117:49]
  assign _T_79 = rawIn_sign ? _T_75 : _T_78; // @[RecFNToIN.scala 114:24]
  assign _T_81 = magGeOne_atOverflowEdge & unroundedInt[30]; // @[RecFNToIN.scala 121:50]
  assign _T_82 = _T_81 & roundCarryBut2; // @[RecFNToIN.scala 122:57]
  assign _T_83 = rawIn_sign | _T_82; // @[RecFNToIN.scala 120:32]
  assign _T_84 = io_signedOut ? _T_79 : _T_83; // @[RecFNToIN.scala 113:20]
  assign _T_85 = _T_71 | _T_84; // @[RecFNToIN.scala 112:40]
  assign _T_87 = ~io_signedOut & rawIn_sign; // @[RecFNToIN.scala 124:28]
  assign _T_88 = _T_87 & roundIncr; // @[RecFNToIN.scala 124:42]
  assign common_overflow = magGeOne ? _T_85 : _T_88; // @[RecFNToIN.scala 111:12]
  assign invalidExc = rawIn_isNaN | rawIn_isInf; // @[RecFNToIN.scala 129:34]
  assign overflow = ~invalidExc & common_overflow; // @[RecFNToIN.scala 130:33]
  assign _T_92 = ~invalidExc & ~common_overflow; // @[RecFNToIN.scala 131:33]
  assign inexact = _T_92 & common_inexact; // @[RecFNToIN.scala 131:54]
  assign _T_100 = {invalidExc,overflow}; // @[Cat.scala 30:58]
  assign io_intExceptionFlags = {_T_100,inexact}; // @[RecFNToIN.scala 142:26]
  assign RecFNToIN_1_covSum = 30'h0;
  assign io_covSum = RecFNToIN_1_covSum;
  assign metaAssert = 1'h0;
endmodule
module INToRecFN(
  input         io_signedIn,
  input  [63:0] io_in,
  input  [2:0]  io_roundingMode,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[INToRecFN.scala 59:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[INToRecFN.scala 59:15]
  wire [7:0] roundAnyRawFNToRecFN_io_in_sExp; // @[INToRecFN.scala 59:15]
  wire [64:0] roundAnyRawFNToRecFN_io_in_sig; // @[INToRecFN.scala 59:15]
  wire [2:0] roundAnyRawFNToRecFN_io_roundingMode; // @[INToRecFN.scala 59:15]
  wire [32:0] roundAnyRawFNToRecFN_io_out; // @[INToRecFN.scala 59:15]
  wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags; // @[INToRecFN.scala 59:15]
  wire [29:0] roundAnyRawFNToRecFN_io_covSum; // @[INToRecFN.scala 59:15]
  wire  roundAnyRawFNToRecFN_metaAssert; // @[INToRecFN.scala 59:15]
  wire  intAsRawFloat_sign; // @[rawFloatFromIN.scala 50:29]
  wire [63:0] _T_14; // @[rawFloatFromIN.scala 51:31]
  wire [63:0] _T_15; // @[rawFloatFromIN.scala 51:24]
  wire [127:0] _T_16; // @[Cat.scala 30:58]
  wire [63:0] _T_21; // @[Bitwise.scala 103:31]
  wire [63:0] _T_23; // @[Bitwise.scala 103:65]
  wire [63:0] _T_25; // @[Bitwise.scala 103:75]
  wire [63:0] _T_26; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_0; // @[Bitwise.scala 103:31]
  wire [63:0] _T_31; // @[Bitwise.scala 103:31]
  wire [63:0] _T_33; // @[Bitwise.scala 103:65]
  wire [63:0] _T_35; // @[Bitwise.scala 103:75]
  wire [63:0] _T_36; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_1; // @[Bitwise.scala 103:31]
  wire [63:0] _T_41; // @[Bitwise.scala 103:31]
  wire [63:0] _T_43; // @[Bitwise.scala 103:65]
  wire [63:0] _T_45; // @[Bitwise.scala 103:75]
  wire [63:0] _T_46; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_2; // @[Bitwise.scala 103:31]
  wire [63:0] _T_51; // @[Bitwise.scala 103:31]
  wire [63:0] _T_53; // @[Bitwise.scala 103:65]
  wire [63:0] _T_55; // @[Bitwise.scala 103:75]
  wire [63:0] _T_56; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_3; // @[Bitwise.scala 103:31]
  wire [63:0] _T_61; // @[Bitwise.scala 103:31]
  wire [63:0] _T_63; // @[Bitwise.scala 103:65]
  wire [63:0] _T_65; // @[Bitwise.scala 103:75]
  wire [63:0] _T_66; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_4; // @[Bitwise.scala 103:31]
  wire [63:0] _T_71; // @[Bitwise.scala 103:31]
  wire [63:0] _T_73; // @[Bitwise.scala 103:65]
  wire [63:0] _T_75; // @[Bitwise.scala 103:75]
  wire [63:0] _T_76; // @[Bitwise.scala 103:39]
  wire [5:0] _T_141; // @[Mux.scala 31:69]
  wire [5:0] _T_142; // @[Mux.scala 31:69]
  wire [5:0] _T_143; // @[Mux.scala 31:69]
  wire [5:0] _T_144; // @[Mux.scala 31:69]
  wire [5:0] _T_145; // @[Mux.scala 31:69]
  wire [5:0] _T_146; // @[Mux.scala 31:69]
  wire [5:0] _T_147; // @[Mux.scala 31:69]
  wire [5:0] _T_148; // @[Mux.scala 31:69]
  wire [5:0] _T_149; // @[Mux.scala 31:69]
  wire [5:0] _T_150; // @[Mux.scala 31:69]
  wire [5:0] _T_151; // @[Mux.scala 31:69]
  wire [5:0] _T_152; // @[Mux.scala 31:69]
  wire [5:0] _T_153; // @[Mux.scala 31:69]
  wire [5:0] _T_154; // @[Mux.scala 31:69]
  wire [5:0] _T_155; // @[Mux.scala 31:69]
  wire [5:0] _T_156; // @[Mux.scala 31:69]
  wire [5:0] _T_157; // @[Mux.scala 31:69]
  wire [5:0] _T_158; // @[Mux.scala 31:69]
  wire [5:0] _T_159; // @[Mux.scala 31:69]
  wire [5:0] _T_160; // @[Mux.scala 31:69]
  wire [5:0] _T_161; // @[Mux.scala 31:69]
  wire [5:0] _T_162; // @[Mux.scala 31:69]
  wire [5:0] _T_163; // @[Mux.scala 31:69]
  wire [5:0] _T_164; // @[Mux.scala 31:69]
  wire [5:0] _T_165; // @[Mux.scala 31:69]
  wire [5:0] _T_166; // @[Mux.scala 31:69]
  wire [5:0] _T_167; // @[Mux.scala 31:69]
  wire [5:0] _T_168; // @[Mux.scala 31:69]
  wire [5:0] _T_169; // @[Mux.scala 31:69]
  wire [5:0] _T_170; // @[Mux.scala 31:69]
  wire [5:0] _T_171; // @[Mux.scala 31:69]
  wire [5:0] _T_172; // @[Mux.scala 31:69]
  wire [5:0] _T_173; // @[Mux.scala 31:69]
  wire [5:0] _T_174; // @[Mux.scala 31:69]
  wire [5:0] _T_175; // @[Mux.scala 31:69]
  wire [5:0] _T_176; // @[Mux.scala 31:69]
  wire [5:0] _T_177; // @[Mux.scala 31:69]
  wire [5:0] _T_178; // @[Mux.scala 31:69]
  wire [5:0] _T_179; // @[Mux.scala 31:69]
  wire [5:0] _T_180; // @[Mux.scala 31:69]
  wire [5:0] _T_181; // @[Mux.scala 31:69]
  wire [5:0] _T_182; // @[Mux.scala 31:69]
  wire [5:0] _T_183; // @[Mux.scala 31:69]
  wire [5:0] _T_184; // @[Mux.scala 31:69]
  wire [5:0] _T_185; // @[Mux.scala 31:69]
  wire [5:0] _T_186; // @[Mux.scala 31:69]
  wire [5:0] _T_187; // @[Mux.scala 31:69]
  wire [5:0] _T_188; // @[Mux.scala 31:69]
  wire [5:0] _T_189; // @[Mux.scala 31:69]
  wire [5:0] _T_190; // @[Mux.scala 31:69]
  wire [5:0] _T_191; // @[Mux.scala 31:69]
  wire [5:0] _T_192; // @[Mux.scala 31:69]
  wire [5:0] _T_193; // @[Mux.scala 31:69]
  wire [5:0] _T_194; // @[Mux.scala 31:69]
  wire [5:0] _T_195; // @[Mux.scala 31:69]
  wire [5:0] _T_196; // @[Mux.scala 31:69]
  wire [5:0] _T_197; // @[Mux.scala 31:69]
  wire [5:0] _T_198; // @[Mux.scala 31:69]
  wire [5:0] _T_199; // @[Mux.scala 31:69]
  wire [5:0] _T_200; // @[Mux.scala 31:69]
  wire [5:0] _T_201; // @[Mux.scala 31:69]
  wire [5:0] _T_202; // @[Mux.scala 31:69]
  wire [5:0] _T_203; // @[Mux.scala 31:69]
  wire [126:0] _GEN_5; // @[rawFloatFromIN.scala 55:22]
  wire [126:0] _T_204; // @[rawFloatFromIN.scala 55:22]
  wire [6:0] _T_211; // @[Cat.scala 30:58]
  wire [29:0] INToRecFN_covSum;
  wire [29:0] roundAnyRawFNToRecFN_sum;
  wire  roundAnyRawFNToRecFN_metaAssert_wire;
  RoundAnyRawFNToRecFN_1 roundAnyRawFNToRecFN ( // @[INToRecFN.scala 59:15]
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),
    .io_out(roundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundAnyRawFNToRecFN_io_covSum),
    .metaAssert(roundAnyRawFNToRecFN_metaAssert)
  );
  assign intAsRawFloat_sign = io_signedIn & io_in[63]; // @[rawFloatFromIN.scala 50:29]
  assign _T_14 = 64'h0 - io_in; // @[rawFloatFromIN.scala 51:31]
  assign _T_15 = intAsRawFloat_sign ? _T_14 : io_in; // @[rawFloatFromIN.scala 51:24]
  assign _T_16 = {64'h0,_T_15}; // @[Cat.scala 30:58]
  assign _T_21 = {{32'd0}, _T_16[63:32]}; // @[Bitwise.scala 103:31]
  assign _T_23 = {_T_16[31:0], 32'h0}; // @[Bitwise.scala 103:65]
  assign _T_25 = _T_23 & 64'hffffffff00000000; // @[Bitwise.scala 103:75]
  assign _T_26 = _T_21 | _T_25; // @[Bitwise.scala 103:39]
  assign _GEN_0 = {{16'd0}, _T_26[63:16]}; // @[Bitwise.scala 103:31]
  assign _T_31 = _GEN_0 & 64'hffff0000ffff; // @[Bitwise.scala 103:31]
  assign _T_33 = {_T_26[47:0], 16'h0}; // @[Bitwise.scala 103:65]
  assign _T_35 = _T_33 & 64'hffff0000ffff0000; // @[Bitwise.scala 103:75]
  assign _T_36 = _T_31 | _T_35; // @[Bitwise.scala 103:39]
  assign _GEN_1 = {{8'd0}, _T_36[63:8]}; // @[Bitwise.scala 103:31]
  assign _T_41 = _GEN_1 & 64'hff00ff00ff00ff; // @[Bitwise.scala 103:31]
  assign _T_43 = {_T_36[55:0], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_45 = _T_43 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 103:75]
  assign _T_46 = _T_41 | _T_45; // @[Bitwise.scala 103:39]
  assign _GEN_2 = {{4'd0}, _T_46[63:4]}; // @[Bitwise.scala 103:31]
  assign _T_51 = _GEN_2 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 103:31]
  assign _T_53 = {_T_46[59:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_55 = _T_53 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 103:75]
  assign _T_56 = _T_51 | _T_55; // @[Bitwise.scala 103:39]
  assign _GEN_3 = {{2'd0}, _T_56[63:2]}; // @[Bitwise.scala 103:31]
  assign _T_61 = _GEN_3 & 64'h3333333333333333; // @[Bitwise.scala 103:31]
  assign _T_63 = {_T_56[61:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_65 = _T_63 & 64'hcccccccccccccccc; // @[Bitwise.scala 103:75]
  assign _T_66 = _T_61 | _T_65; // @[Bitwise.scala 103:39]
  assign _GEN_4 = {{1'd0}, _T_66[63:1]}; // @[Bitwise.scala 103:31]
  assign _T_71 = _GEN_4 & 64'h5555555555555555; // @[Bitwise.scala 103:31]
  assign _T_73 = {_T_66[62:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_75 = _T_73 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 103:75]
  assign _T_76 = _T_71 | _T_75; // @[Bitwise.scala 103:39]
  assign _T_141 = _T_76[62] ? 6'h3e : 6'h3f; // @[Mux.scala 31:69]
  assign _T_142 = _T_76[61] ? 6'h3d : _T_141; // @[Mux.scala 31:69]
  assign _T_143 = _T_76[60] ? 6'h3c : _T_142; // @[Mux.scala 31:69]
  assign _T_144 = _T_76[59] ? 6'h3b : _T_143; // @[Mux.scala 31:69]
  assign _T_145 = _T_76[58] ? 6'h3a : _T_144; // @[Mux.scala 31:69]
  assign _T_146 = _T_76[57] ? 6'h39 : _T_145; // @[Mux.scala 31:69]
  assign _T_147 = _T_76[56] ? 6'h38 : _T_146; // @[Mux.scala 31:69]
  assign _T_148 = _T_76[55] ? 6'h37 : _T_147; // @[Mux.scala 31:69]
  assign _T_149 = _T_76[54] ? 6'h36 : _T_148; // @[Mux.scala 31:69]
  assign _T_150 = _T_76[53] ? 6'h35 : _T_149; // @[Mux.scala 31:69]
  assign _T_151 = _T_76[52] ? 6'h34 : _T_150; // @[Mux.scala 31:69]
  assign _T_152 = _T_76[51] ? 6'h33 : _T_151; // @[Mux.scala 31:69]
  assign _T_153 = _T_76[50] ? 6'h32 : _T_152; // @[Mux.scala 31:69]
  assign _T_154 = _T_76[49] ? 6'h31 : _T_153; // @[Mux.scala 31:69]
  assign _T_155 = _T_76[48] ? 6'h30 : _T_154; // @[Mux.scala 31:69]
  assign _T_156 = _T_76[47] ? 6'h2f : _T_155; // @[Mux.scala 31:69]
  assign _T_157 = _T_76[46] ? 6'h2e : _T_156; // @[Mux.scala 31:69]
  assign _T_158 = _T_76[45] ? 6'h2d : _T_157; // @[Mux.scala 31:69]
  assign _T_159 = _T_76[44] ? 6'h2c : _T_158; // @[Mux.scala 31:69]
  assign _T_160 = _T_76[43] ? 6'h2b : _T_159; // @[Mux.scala 31:69]
  assign _T_161 = _T_76[42] ? 6'h2a : _T_160; // @[Mux.scala 31:69]
  assign _T_162 = _T_76[41] ? 6'h29 : _T_161; // @[Mux.scala 31:69]
  assign _T_163 = _T_76[40] ? 6'h28 : _T_162; // @[Mux.scala 31:69]
  assign _T_164 = _T_76[39] ? 6'h27 : _T_163; // @[Mux.scala 31:69]
  assign _T_165 = _T_76[38] ? 6'h26 : _T_164; // @[Mux.scala 31:69]
  assign _T_166 = _T_76[37] ? 6'h25 : _T_165; // @[Mux.scala 31:69]
  assign _T_167 = _T_76[36] ? 6'h24 : _T_166; // @[Mux.scala 31:69]
  assign _T_168 = _T_76[35] ? 6'h23 : _T_167; // @[Mux.scala 31:69]
  assign _T_169 = _T_76[34] ? 6'h22 : _T_168; // @[Mux.scala 31:69]
  assign _T_170 = _T_76[33] ? 6'h21 : _T_169; // @[Mux.scala 31:69]
  assign _T_171 = _T_76[32] ? 6'h20 : _T_170; // @[Mux.scala 31:69]
  assign _T_172 = _T_76[31] ? 6'h1f : _T_171; // @[Mux.scala 31:69]
  assign _T_173 = _T_76[30] ? 6'h1e : _T_172; // @[Mux.scala 31:69]
  assign _T_174 = _T_76[29] ? 6'h1d : _T_173; // @[Mux.scala 31:69]
  assign _T_175 = _T_76[28] ? 6'h1c : _T_174; // @[Mux.scala 31:69]
  assign _T_176 = _T_76[27] ? 6'h1b : _T_175; // @[Mux.scala 31:69]
  assign _T_177 = _T_76[26] ? 6'h1a : _T_176; // @[Mux.scala 31:69]
  assign _T_178 = _T_76[25] ? 6'h19 : _T_177; // @[Mux.scala 31:69]
  assign _T_179 = _T_76[24] ? 6'h18 : _T_178; // @[Mux.scala 31:69]
  assign _T_180 = _T_76[23] ? 6'h17 : _T_179; // @[Mux.scala 31:69]
  assign _T_181 = _T_76[22] ? 6'h16 : _T_180; // @[Mux.scala 31:69]
  assign _T_182 = _T_76[21] ? 6'h15 : _T_181; // @[Mux.scala 31:69]
  assign _T_183 = _T_76[20] ? 6'h14 : _T_182; // @[Mux.scala 31:69]
  assign _T_184 = _T_76[19] ? 6'h13 : _T_183; // @[Mux.scala 31:69]
  assign _T_185 = _T_76[18] ? 6'h12 : _T_184; // @[Mux.scala 31:69]
  assign _T_186 = _T_76[17] ? 6'h11 : _T_185; // @[Mux.scala 31:69]
  assign _T_187 = _T_76[16] ? 6'h10 : _T_186; // @[Mux.scala 31:69]
  assign _T_188 = _T_76[15] ? 6'hf : _T_187; // @[Mux.scala 31:69]
  assign _T_189 = _T_76[14] ? 6'he : _T_188; // @[Mux.scala 31:69]
  assign _T_190 = _T_76[13] ? 6'hd : _T_189; // @[Mux.scala 31:69]
  assign _T_191 = _T_76[12] ? 6'hc : _T_190; // @[Mux.scala 31:69]
  assign _T_192 = _T_76[11] ? 6'hb : _T_191; // @[Mux.scala 31:69]
  assign _T_193 = _T_76[10] ? 6'ha : _T_192; // @[Mux.scala 31:69]
  assign _T_194 = _T_76[9] ? 6'h9 : _T_193; // @[Mux.scala 31:69]
  assign _T_195 = _T_76[8] ? 6'h8 : _T_194; // @[Mux.scala 31:69]
  assign _T_196 = _T_76[7] ? 6'h7 : _T_195; // @[Mux.scala 31:69]
  assign _T_197 = _T_76[6] ? 6'h6 : _T_196; // @[Mux.scala 31:69]
  assign _T_198 = _T_76[5] ? 6'h5 : _T_197; // @[Mux.scala 31:69]
  assign _T_199 = _T_76[4] ? 6'h4 : _T_198; // @[Mux.scala 31:69]
  assign _T_200 = _T_76[3] ? 6'h3 : _T_199; // @[Mux.scala 31:69]
  assign _T_201 = _T_76[2] ? 6'h2 : _T_200; // @[Mux.scala 31:69]
  assign _T_202 = _T_76[1] ? 6'h1 : _T_201; // @[Mux.scala 31:69]
  assign _T_203 = _T_76[0] ? 6'h0 : _T_202; // @[Mux.scala 31:69]
  assign _GEN_5 = {{63'd0}, _T_16[63:0]}; // @[rawFloatFromIN.scala 55:22]
  assign _T_204 = _GEN_5 << _T_203; // @[rawFloatFromIN.scala 55:22]
  assign _T_211 = {1'h1,~_T_203}; // @[Cat.scala 30:58]
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[INToRecFN.scala 72:23]
  assign io_exceptionFlags = roundAnyRawFNToRecFN_io_exceptionFlags; // @[INToRecFN.scala 73:23]
  assign roundAnyRawFNToRecFN_io_in_isZero = ~_T_204[63]; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_signedIn & io_in[63]; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = {1'b0,$signed(_T_211)}; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sig = {{1'd0}, _T_204[63:0]}; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[INToRecFN.scala 70:44]
  assign INToRecFN_covSum = 30'h0;
  assign roundAnyRawFNToRecFN_sum = INToRecFN_covSum + roundAnyRawFNToRecFN_io_covSum;
  assign io_covSum = roundAnyRawFNToRecFN_sum;
  assign roundAnyRawFNToRecFN_metaAssert_wire = roundAnyRawFNToRecFN_metaAssert;
  assign metaAssert = roundAnyRawFNToRecFN_metaAssert_wire;
endmodule
module INToRecFN_1(
  input         io_signedIn,
  input  [63:0] io_in,
  input  [2:0]  io_roundingMode,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[INToRecFN.scala 59:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[INToRecFN.scala 59:15]
  wire [7:0] roundAnyRawFNToRecFN_io_in_sExp; // @[INToRecFN.scala 59:15]
  wire [64:0] roundAnyRawFNToRecFN_io_in_sig; // @[INToRecFN.scala 59:15]
  wire [2:0] roundAnyRawFNToRecFN_io_roundingMode; // @[INToRecFN.scala 59:15]
  wire [64:0] roundAnyRawFNToRecFN_io_out; // @[INToRecFN.scala 59:15]
  wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags; // @[INToRecFN.scala 59:15]
  wire [29:0] roundAnyRawFNToRecFN_io_covSum; // @[INToRecFN.scala 59:15]
  wire  roundAnyRawFNToRecFN_metaAssert; // @[INToRecFN.scala 59:15]
  wire  intAsRawFloat_sign; // @[rawFloatFromIN.scala 50:29]
  wire [63:0] _T_14; // @[rawFloatFromIN.scala 51:31]
  wire [63:0] _T_15; // @[rawFloatFromIN.scala 51:24]
  wire [127:0] _T_16; // @[Cat.scala 30:58]
  wire [63:0] _T_21; // @[Bitwise.scala 103:31]
  wire [63:0] _T_23; // @[Bitwise.scala 103:65]
  wire [63:0] _T_25; // @[Bitwise.scala 103:75]
  wire [63:0] _T_26; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_0; // @[Bitwise.scala 103:31]
  wire [63:0] _T_31; // @[Bitwise.scala 103:31]
  wire [63:0] _T_33; // @[Bitwise.scala 103:65]
  wire [63:0] _T_35; // @[Bitwise.scala 103:75]
  wire [63:0] _T_36; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_1; // @[Bitwise.scala 103:31]
  wire [63:0] _T_41; // @[Bitwise.scala 103:31]
  wire [63:0] _T_43; // @[Bitwise.scala 103:65]
  wire [63:0] _T_45; // @[Bitwise.scala 103:75]
  wire [63:0] _T_46; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_2; // @[Bitwise.scala 103:31]
  wire [63:0] _T_51; // @[Bitwise.scala 103:31]
  wire [63:0] _T_53; // @[Bitwise.scala 103:65]
  wire [63:0] _T_55; // @[Bitwise.scala 103:75]
  wire [63:0] _T_56; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_3; // @[Bitwise.scala 103:31]
  wire [63:0] _T_61; // @[Bitwise.scala 103:31]
  wire [63:0] _T_63; // @[Bitwise.scala 103:65]
  wire [63:0] _T_65; // @[Bitwise.scala 103:75]
  wire [63:0] _T_66; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_4; // @[Bitwise.scala 103:31]
  wire [63:0] _T_71; // @[Bitwise.scala 103:31]
  wire [63:0] _T_73; // @[Bitwise.scala 103:65]
  wire [63:0] _T_75; // @[Bitwise.scala 103:75]
  wire [63:0] _T_76; // @[Bitwise.scala 103:39]
  wire [5:0] _T_141; // @[Mux.scala 31:69]
  wire [5:0] _T_142; // @[Mux.scala 31:69]
  wire [5:0] _T_143; // @[Mux.scala 31:69]
  wire [5:0] _T_144; // @[Mux.scala 31:69]
  wire [5:0] _T_145; // @[Mux.scala 31:69]
  wire [5:0] _T_146; // @[Mux.scala 31:69]
  wire [5:0] _T_147; // @[Mux.scala 31:69]
  wire [5:0] _T_148; // @[Mux.scala 31:69]
  wire [5:0] _T_149; // @[Mux.scala 31:69]
  wire [5:0] _T_150; // @[Mux.scala 31:69]
  wire [5:0] _T_151; // @[Mux.scala 31:69]
  wire [5:0] _T_152; // @[Mux.scala 31:69]
  wire [5:0] _T_153; // @[Mux.scala 31:69]
  wire [5:0] _T_154; // @[Mux.scala 31:69]
  wire [5:0] _T_155; // @[Mux.scala 31:69]
  wire [5:0] _T_156; // @[Mux.scala 31:69]
  wire [5:0] _T_157; // @[Mux.scala 31:69]
  wire [5:0] _T_158; // @[Mux.scala 31:69]
  wire [5:0] _T_159; // @[Mux.scala 31:69]
  wire [5:0] _T_160; // @[Mux.scala 31:69]
  wire [5:0] _T_161; // @[Mux.scala 31:69]
  wire [5:0] _T_162; // @[Mux.scala 31:69]
  wire [5:0] _T_163; // @[Mux.scala 31:69]
  wire [5:0] _T_164; // @[Mux.scala 31:69]
  wire [5:0] _T_165; // @[Mux.scala 31:69]
  wire [5:0] _T_166; // @[Mux.scala 31:69]
  wire [5:0] _T_167; // @[Mux.scala 31:69]
  wire [5:0] _T_168; // @[Mux.scala 31:69]
  wire [5:0] _T_169; // @[Mux.scala 31:69]
  wire [5:0] _T_170; // @[Mux.scala 31:69]
  wire [5:0] _T_171; // @[Mux.scala 31:69]
  wire [5:0] _T_172; // @[Mux.scala 31:69]
  wire [5:0] _T_173; // @[Mux.scala 31:69]
  wire [5:0] _T_174; // @[Mux.scala 31:69]
  wire [5:0] _T_175; // @[Mux.scala 31:69]
  wire [5:0] _T_176; // @[Mux.scala 31:69]
  wire [5:0] _T_177; // @[Mux.scala 31:69]
  wire [5:0] _T_178; // @[Mux.scala 31:69]
  wire [5:0] _T_179; // @[Mux.scala 31:69]
  wire [5:0] _T_180; // @[Mux.scala 31:69]
  wire [5:0] _T_181; // @[Mux.scala 31:69]
  wire [5:0] _T_182; // @[Mux.scala 31:69]
  wire [5:0] _T_183; // @[Mux.scala 31:69]
  wire [5:0] _T_184; // @[Mux.scala 31:69]
  wire [5:0] _T_185; // @[Mux.scala 31:69]
  wire [5:0] _T_186; // @[Mux.scala 31:69]
  wire [5:0] _T_187; // @[Mux.scala 31:69]
  wire [5:0] _T_188; // @[Mux.scala 31:69]
  wire [5:0] _T_189; // @[Mux.scala 31:69]
  wire [5:0] _T_190; // @[Mux.scala 31:69]
  wire [5:0] _T_191; // @[Mux.scala 31:69]
  wire [5:0] _T_192; // @[Mux.scala 31:69]
  wire [5:0] _T_193; // @[Mux.scala 31:69]
  wire [5:0] _T_194; // @[Mux.scala 31:69]
  wire [5:0] _T_195; // @[Mux.scala 31:69]
  wire [5:0] _T_196; // @[Mux.scala 31:69]
  wire [5:0] _T_197; // @[Mux.scala 31:69]
  wire [5:0] _T_198; // @[Mux.scala 31:69]
  wire [5:0] _T_199; // @[Mux.scala 31:69]
  wire [5:0] _T_200; // @[Mux.scala 31:69]
  wire [5:0] _T_201; // @[Mux.scala 31:69]
  wire [5:0] _T_202; // @[Mux.scala 31:69]
  wire [5:0] _T_203; // @[Mux.scala 31:69]
  wire [126:0] _GEN_5; // @[rawFloatFromIN.scala 55:22]
  wire [126:0] _T_204; // @[rawFloatFromIN.scala 55:22]
  wire [6:0] _T_211; // @[Cat.scala 30:58]
  wire [29:0] INToRecFN_1_covSum;
  wire [29:0] roundAnyRawFNToRecFN_sum;
  wire  roundAnyRawFNToRecFN_metaAssert_wire;
  RoundAnyRawFNToRecFN_2 roundAnyRawFNToRecFN ( // @[INToRecFN.scala 59:15]
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),
    .io_out(roundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundAnyRawFNToRecFN_io_covSum),
    .metaAssert(roundAnyRawFNToRecFN_metaAssert)
  );
  assign intAsRawFloat_sign = io_signedIn & io_in[63]; // @[rawFloatFromIN.scala 50:29]
  assign _T_14 = 64'h0 - io_in; // @[rawFloatFromIN.scala 51:31]
  assign _T_15 = intAsRawFloat_sign ? _T_14 : io_in; // @[rawFloatFromIN.scala 51:24]
  assign _T_16 = {64'h0,_T_15}; // @[Cat.scala 30:58]
  assign _T_21 = {{32'd0}, _T_16[63:32]}; // @[Bitwise.scala 103:31]
  assign _T_23 = {_T_16[31:0], 32'h0}; // @[Bitwise.scala 103:65]
  assign _T_25 = _T_23 & 64'hffffffff00000000; // @[Bitwise.scala 103:75]
  assign _T_26 = _T_21 | _T_25; // @[Bitwise.scala 103:39]
  assign _GEN_0 = {{16'd0}, _T_26[63:16]}; // @[Bitwise.scala 103:31]
  assign _T_31 = _GEN_0 & 64'hffff0000ffff; // @[Bitwise.scala 103:31]
  assign _T_33 = {_T_26[47:0], 16'h0}; // @[Bitwise.scala 103:65]
  assign _T_35 = _T_33 & 64'hffff0000ffff0000; // @[Bitwise.scala 103:75]
  assign _T_36 = _T_31 | _T_35; // @[Bitwise.scala 103:39]
  assign _GEN_1 = {{8'd0}, _T_36[63:8]}; // @[Bitwise.scala 103:31]
  assign _T_41 = _GEN_1 & 64'hff00ff00ff00ff; // @[Bitwise.scala 103:31]
  assign _T_43 = {_T_36[55:0], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_45 = _T_43 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 103:75]
  assign _T_46 = _T_41 | _T_45; // @[Bitwise.scala 103:39]
  assign _GEN_2 = {{4'd0}, _T_46[63:4]}; // @[Bitwise.scala 103:31]
  assign _T_51 = _GEN_2 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 103:31]
  assign _T_53 = {_T_46[59:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_55 = _T_53 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 103:75]
  assign _T_56 = _T_51 | _T_55; // @[Bitwise.scala 103:39]
  assign _GEN_3 = {{2'd0}, _T_56[63:2]}; // @[Bitwise.scala 103:31]
  assign _T_61 = _GEN_3 & 64'h3333333333333333; // @[Bitwise.scala 103:31]
  assign _T_63 = {_T_56[61:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_65 = _T_63 & 64'hcccccccccccccccc; // @[Bitwise.scala 103:75]
  assign _T_66 = _T_61 | _T_65; // @[Bitwise.scala 103:39]
  assign _GEN_4 = {{1'd0}, _T_66[63:1]}; // @[Bitwise.scala 103:31]
  assign _T_71 = _GEN_4 & 64'h5555555555555555; // @[Bitwise.scala 103:31]
  assign _T_73 = {_T_66[62:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_75 = _T_73 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 103:75]
  assign _T_76 = _T_71 | _T_75; // @[Bitwise.scala 103:39]
  assign _T_141 = _T_76[62] ? 6'h3e : 6'h3f; // @[Mux.scala 31:69]
  assign _T_142 = _T_76[61] ? 6'h3d : _T_141; // @[Mux.scala 31:69]
  assign _T_143 = _T_76[60] ? 6'h3c : _T_142; // @[Mux.scala 31:69]
  assign _T_144 = _T_76[59] ? 6'h3b : _T_143; // @[Mux.scala 31:69]
  assign _T_145 = _T_76[58] ? 6'h3a : _T_144; // @[Mux.scala 31:69]
  assign _T_146 = _T_76[57] ? 6'h39 : _T_145; // @[Mux.scala 31:69]
  assign _T_147 = _T_76[56] ? 6'h38 : _T_146; // @[Mux.scala 31:69]
  assign _T_148 = _T_76[55] ? 6'h37 : _T_147; // @[Mux.scala 31:69]
  assign _T_149 = _T_76[54] ? 6'h36 : _T_148; // @[Mux.scala 31:69]
  assign _T_150 = _T_76[53] ? 6'h35 : _T_149; // @[Mux.scala 31:69]
  assign _T_151 = _T_76[52] ? 6'h34 : _T_150; // @[Mux.scala 31:69]
  assign _T_152 = _T_76[51] ? 6'h33 : _T_151; // @[Mux.scala 31:69]
  assign _T_153 = _T_76[50] ? 6'h32 : _T_152; // @[Mux.scala 31:69]
  assign _T_154 = _T_76[49] ? 6'h31 : _T_153; // @[Mux.scala 31:69]
  assign _T_155 = _T_76[48] ? 6'h30 : _T_154; // @[Mux.scala 31:69]
  assign _T_156 = _T_76[47] ? 6'h2f : _T_155; // @[Mux.scala 31:69]
  assign _T_157 = _T_76[46] ? 6'h2e : _T_156; // @[Mux.scala 31:69]
  assign _T_158 = _T_76[45] ? 6'h2d : _T_157; // @[Mux.scala 31:69]
  assign _T_159 = _T_76[44] ? 6'h2c : _T_158; // @[Mux.scala 31:69]
  assign _T_160 = _T_76[43] ? 6'h2b : _T_159; // @[Mux.scala 31:69]
  assign _T_161 = _T_76[42] ? 6'h2a : _T_160; // @[Mux.scala 31:69]
  assign _T_162 = _T_76[41] ? 6'h29 : _T_161; // @[Mux.scala 31:69]
  assign _T_163 = _T_76[40] ? 6'h28 : _T_162; // @[Mux.scala 31:69]
  assign _T_164 = _T_76[39] ? 6'h27 : _T_163; // @[Mux.scala 31:69]
  assign _T_165 = _T_76[38] ? 6'h26 : _T_164; // @[Mux.scala 31:69]
  assign _T_166 = _T_76[37] ? 6'h25 : _T_165; // @[Mux.scala 31:69]
  assign _T_167 = _T_76[36] ? 6'h24 : _T_166; // @[Mux.scala 31:69]
  assign _T_168 = _T_76[35] ? 6'h23 : _T_167; // @[Mux.scala 31:69]
  assign _T_169 = _T_76[34] ? 6'h22 : _T_168; // @[Mux.scala 31:69]
  assign _T_170 = _T_76[33] ? 6'h21 : _T_169; // @[Mux.scala 31:69]
  assign _T_171 = _T_76[32] ? 6'h20 : _T_170; // @[Mux.scala 31:69]
  assign _T_172 = _T_76[31] ? 6'h1f : _T_171; // @[Mux.scala 31:69]
  assign _T_173 = _T_76[30] ? 6'h1e : _T_172; // @[Mux.scala 31:69]
  assign _T_174 = _T_76[29] ? 6'h1d : _T_173; // @[Mux.scala 31:69]
  assign _T_175 = _T_76[28] ? 6'h1c : _T_174; // @[Mux.scala 31:69]
  assign _T_176 = _T_76[27] ? 6'h1b : _T_175; // @[Mux.scala 31:69]
  assign _T_177 = _T_76[26] ? 6'h1a : _T_176; // @[Mux.scala 31:69]
  assign _T_178 = _T_76[25] ? 6'h19 : _T_177; // @[Mux.scala 31:69]
  assign _T_179 = _T_76[24] ? 6'h18 : _T_178; // @[Mux.scala 31:69]
  assign _T_180 = _T_76[23] ? 6'h17 : _T_179; // @[Mux.scala 31:69]
  assign _T_181 = _T_76[22] ? 6'h16 : _T_180; // @[Mux.scala 31:69]
  assign _T_182 = _T_76[21] ? 6'h15 : _T_181; // @[Mux.scala 31:69]
  assign _T_183 = _T_76[20] ? 6'h14 : _T_182; // @[Mux.scala 31:69]
  assign _T_184 = _T_76[19] ? 6'h13 : _T_183; // @[Mux.scala 31:69]
  assign _T_185 = _T_76[18] ? 6'h12 : _T_184; // @[Mux.scala 31:69]
  assign _T_186 = _T_76[17] ? 6'h11 : _T_185; // @[Mux.scala 31:69]
  assign _T_187 = _T_76[16] ? 6'h10 : _T_186; // @[Mux.scala 31:69]
  assign _T_188 = _T_76[15] ? 6'hf : _T_187; // @[Mux.scala 31:69]
  assign _T_189 = _T_76[14] ? 6'he : _T_188; // @[Mux.scala 31:69]
  assign _T_190 = _T_76[13] ? 6'hd : _T_189; // @[Mux.scala 31:69]
  assign _T_191 = _T_76[12] ? 6'hc : _T_190; // @[Mux.scala 31:69]
  assign _T_192 = _T_76[11] ? 6'hb : _T_191; // @[Mux.scala 31:69]
  assign _T_193 = _T_76[10] ? 6'ha : _T_192; // @[Mux.scala 31:69]
  assign _T_194 = _T_76[9] ? 6'h9 : _T_193; // @[Mux.scala 31:69]
  assign _T_195 = _T_76[8] ? 6'h8 : _T_194; // @[Mux.scala 31:69]
  assign _T_196 = _T_76[7] ? 6'h7 : _T_195; // @[Mux.scala 31:69]
  assign _T_197 = _T_76[6] ? 6'h6 : _T_196; // @[Mux.scala 31:69]
  assign _T_198 = _T_76[5] ? 6'h5 : _T_197; // @[Mux.scala 31:69]
  assign _T_199 = _T_76[4] ? 6'h4 : _T_198; // @[Mux.scala 31:69]
  assign _T_200 = _T_76[3] ? 6'h3 : _T_199; // @[Mux.scala 31:69]
  assign _T_201 = _T_76[2] ? 6'h2 : _T_200; // @[Mux.scala 31:69]
  assign _T_202 = _T_76[1] ? 6'h1 : _T_201; // @[Mux.scala 31:69]
  assign _T_203 = _T_76[0] ? 6'h0 : _T_202; // @[Mux.scala 31:69]
  assign _GEN_5 = {{63'd0}, _T_16[63:0]}; // @[rawFloatFromIN.scala 55:22]
  assign _T_204 = _GEN_5 << _T_203; // @[rawFloatFromIN.scala 55:22]
  assign _T_211 = {1'h1,~_T_203}; // @[Cat.scala 30:58]
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[INToRecFN.scala 72:23]
  assign io_exceptionFlags = roundAnyRawFNToRecFN_io_exceptionFlags; // @[INToRecFN.scala 73:23]
  assign roundAnyRawFNToRecFN_io_in_isZero = ~_T_204[63]; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_signedIn & io_in[63]; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = {1'b0,$signed(_T_211)}; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sig = {{1'd0}, _T_204[63:0]}; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[INToRecFN.scala 70:44]
  assign INToRecFN_1_covSum = 30'h0;
  assign roundAnyRawFNToRecFN_sum = INToRecFN_1_covSum + roundAnyRawFNToRecFN_io_covSum;
  assign io_covSum = roundAnyRawFNToRecFN_sum;
  assign roundAnyRawFNToRecFN_metaAssert_wire = roundAnyRawFNToRecFN_metaAssert;
  assign metaAssert = roundAnyRawFNToRecFN_metaAssert_wire;
endmodule
module RecFNToRecFN(
  input  [64:0] io_in,
  input  [2:0]  io_roundingMode,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  RoundAnyRawFNToRecFN_io_invalidExc; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_io_in_isNaN; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_io_in_isInf; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_io_in_isZero; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_io_in_sign; // @[RecFNToRecFN.scala 72:19]
  wire [12:0] RoundAnyRawFNToRecFN_io_in_sExp; // @[RecFNToRecFN.scala 72:19]
  wire [53:0] RoundAnyRawFNToRecFN_io_in_sig; // @[RecFNToRecFN.scala 72:19]
  wire [2:0] RoundAnyRawFNToRecFN_io_roundingMode; // @[RecFNToRecFN.scala 72:19]
  wire [32:0] RoundAnyRawFNToRecFN_io_out; // @[RecFNToRecFN.scala 72:19]
  wire [4:0] RoundAnyRawFNToRecFN_io_exceptionFlags; // @[RecFNToRecFN.scala 72:19]
  wire [29:0] RoundAnyRawFNToRecFN_io_covSum; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_metaAssert; // @[RecFNToRecFN.scala 72:19]
  wire  rawIn_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_13; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawIn_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire [1:0] _T_24; // @[Cat.scala 30:58]
  wire [53:0] rawIn_sig; // @[Cat.scala 30:58]
  wire [29:0] RecFNToRecFN_covSum;
  wire [29:0] RoundAnyRawFNToRecFN_sum;
  wire  RoundAnyRawFNToRecFN_metaAssert_wire;
  RoundAnyRawFNToRecFN_3 RoundAnyRawFNToRecFN ( // @[RecFNToRecFN.scala 72:19]
    .io_invalidExc(RoundAnyRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(RoundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(RoundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(RoundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(RoundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(RoundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(RoundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(RoundAnyRawFNToRecFN_io_roundingMode),
    .io_out(RoundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(RoundAnyRawFNToRecFN_io_exceptionFlags),
    .io_covSum(RoundAnyRawFNToRecFN_io_covSum),
    .metaAssert(RoundAnyRawFNToRecFN_metaAssert)
  );
  assign rawIn_isZero = io_in[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_13 = io_in[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawIn_isNaN = _T_13 & io_in[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign _T_24 = {1'h0,~rawIn_isZero}; // @[Cat.scala 30:58]
  assign rawIn_sig = {1'h0,~rawIn_isZero,io_in[51:0]}; // @[Cat.scala 30:58]
  assign io_out = RoundAnyRawFNToRecFN_io_out; // @[RecFNToRecFN.scala 85:27]
  assign io_exceptionFlags = RoundAnyRawFNToRecFN_io_exceptionFlags; // @[RecFNToRecFN.scala 86:27]
  assign RoundAnyRawFNToRecFN_io_invalidExc = rawIn_isNaN & ~rawIn_sig[51]; // @[RecFNToRecFN.scala 80:48]
  assign RoundAnyRawFNToRecFN_io_in_isNaN = _T_13 & io_in[61]; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_isInf = _T_13 & ~io_in[61]; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_isZero = io_in[63:61] == 3'h0; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_sign = io_in[64]; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_sExp = {1'b0,$signed(io_in[63:52])}; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_sig = {_T_24,io_in[51:0]}; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[RecFNToRecFN.scala 83:48]
  assign RecFNToRecFN_covSum = 30'h0;
  assign RoundAnyRawFNToRecFN_sum = RecFNToRecFN_covSum + RoundAnyRawFNToRecFN_io_covSum;
  assign io_covSum = RoundAnyRawFNToRecFN_sum;
  assign RoundAnyRawFNToRecFN_metaAssert_wire = RoundAnyRawFNToRecFN_metaAssert;
  assign metaAssert = RoundAnyRawFNToRecFN_metaAssert_wire;
endmodule
module MulAddRecFNPipe_1(
  input         clock,
  input         reset,
  input         io_validin,
  input  [1:0]  io_op,
  input  [64:0] io_a,
  input  [64:0] io_b,
  input  [64:0] io_c,
  input  [2:0]  io_roundingMode,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags,
  output        io_validout,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [1:0] mulAddRecFNToRaw_preMul_io_op; // @[FPU.scala 580:15]
  wire [64:0] mulAddRecFNToRaw_preMul_io_a; // @[FPU.scala 580:15]
  wire [64:0] mulAddRecFNToRaw_preMul_io_b; // @[FPU.scala 580:15]
  wire [64:0] mulAddRecFNToRaw_preMul_io_c; // @[FPU.scala 580:15]
  wire [52:0] mulAddRecFNToRaw_preMul_io_mulAddA; // @[FPU.scala 580:15]
  wire [52:0] mulAddRecFNToRaw_preMul_io_mulAddB; // @[FPU.scala 580:15]
  wire [105:0] mulAddRecFNToRaw_preMul_io_mulAddC; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[FPU.scala 580:15]
  wire [12:0] mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[FPU.scala 580:15]
  wire [5:0] mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[FPU.scala 580:15]
  wire [54:0] mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[FPU.scala 580:15]
  wire [29:0] mulAddRecFNToRaw_preMul_io_covSum; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_preMul_metaAssert; // @[FPU.scala 580:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_signProd; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC; // @[FPU.scala 582:15]
  wire [12:0] mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant; // @[FPU.scala 582:15]
  wire [5:0] mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist; // @[FPU.scala 582:15]
  wire [54:0] mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC; // @[FPU.scala 582:15]
  wire [106:0] mulAddRecFNToRaw_postMul_io_mulAddResult; // @[FPU.scala 582:15]
  wire [2:0] mulAddRecFNToRaw_postMul_io_roundingMode; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_invalidExc; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[FPU.scala 582:15]
  wire [12:0] mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[FPU.scala 582:15]
  wire [55:0] mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[FPU.scala 582:15]
  wire [29:0] mulAddRecFNToRaw_postMul_io_covSum; // @[FPU.scala 582:15]
  wire  mulAddRecFNToRaw_postMul_metaAssert; // @[FPU.scala 582:15]
  wire  roundRawFNToRecFN_io_invalidExc; // @[FPU.scala 608:35]
  wire  roundRawFNToRecFN_io_infiniteExc; // @[FPU.scala 608:35]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[FPU.scala 608:35]
  wire  roundRawFNToRecFN_io_in_isInf; // @[FPU.scala 608:35]
  wire  roundRawFNToRecFN_io_in_isZero; // @[FPU.scala 608:35]
  wire  roundRawFNToRecFN_io_in_sign; // @[FPU.scala 608:35]
  wire [12:0] roundRawFNToRecFN_io_in_sExp; // @[FPU.scala 608:35]
  wire [55:0] roundRawFNToRecFN_io_in_sig; // @[FPU.scala 608:35]
  wire [2:0] roundRawFNToRecFN_io_roundingMode; // @[FPU.scala 608:35]
  wire  roundRawFNToRecFN_io_detectTininess; // @[FPU.scala 608:35]
  wire [64:0] roundRawFNToRecFN_io_out; // @[FPU.scala 608:35]
  wire [4:0] roundRawFNToRecFN_io_exceptionFlags; // @[FPU.scala 608:35]
  wire [29:0] roundRawFNToRecFN_io_covSum; // @[FPU.scala 608:35]
  wire  roundRawFNToRecFN_metaAssert; // @[FPU.scala 608:35]
  wire [105:0] _T_14; // @[FPU.scala 590:45]
  wire [106:0] mulAddResult; // @[FPU.scala 591:50]
  reg  _T_21_isSigNaNAny; // @[Reg.scala 11:16]
  reg [31:0] _RAND_0;
  reg  _T_21_isNaNAOrB; // @[Reg.scala 11:16]
  reg [31:0] _RAND_1;
  reg  _T_21_isInfA; // @[Reg.scala 11:16]
  reg [31:0] _RAND_2;
  reg  _T_21_isZeroA; // @[Reg.scala 11:16]
  reg [31:0] _RAND_3;
  reg  _T_21_isInfB; // @[Reg.scala 11:16]
  reg [31:0] _RAND_4;
  reg  _T_21_isZeroB; // @[Reg.scala 11:16]
  reg [31:0] _RAND_5;
  reg  _T_21_signProd; // @[Reg.scala 11:16]
  reg [31:0] _RAND_6;
  reg  _T_21_isNaNC; // @[Reg.scala 11:16]
  reg [31:0] _RAND_7;
  reg  _T_21_isInfC; // @[Reg.scala 11:16]
  reg [31:0] _RAND_8;
  reg  _T_21_isZeroC; // @[Reg.scala 11:16]
  reg [31:0] _RAND_9;
  reg [12:0] _T_21_sExpSum; // @[Reg.scala 11:16]
  reg [31:0] _RAND_10;
  reg  _T_21_doSubMags; // @[Reg.scala 11:16]
  reg [31:0] _RAND_11;
  reg  _T_21_CIsDominant; // @[Reg.scala 11:16]
  reg [31:0] _RAND_12;
  reg [5:0] _T_21_CDom_CAlignDist; // @[Reg.scala 11:16]
  reg [31:0] _RAND_13;
  reg [54:0] _T_21_highAlignedSigC; // @[Reg.scala 11:16]
  reg [63:0] _RAND_14;
  reg  _T_21_bit0AlignedSigC; // @[Reg.scala 11:16]
  reg [31:0] _RAND_15;
  reg [106:0] _T_30; // @[Reg.scala 11:16]
  reg [127:0] _RAND_16;
  reg [2:0] _T_39; // @[Reg.scala 11:16]
  reg [31:0] _RAND_17;
  reg [2:0] roundingMode_stage0; // @[Reg.scala 11:16]
  reg [31:0] _RAND_18;
  reg  detectTininess_stage0; // @[Reg.scala 11:16]
  reg [31:0] _RAND_19;
  reg  valid_stage0; // @[Valid.scala 48:22]
  reg [31:0] _RAND_20;
  reg  _T_75; // @[Reg.scala 11:16]
  reg [31:0] _RAND_21;
  reg  _T_84_isNaN; // @[Reg.scala 11:16]
  reg [31:0] _RAND_22;
  reg  _T_84_isInf; // @[Reg.scala 11:16]
  reg [31:0] _RAND_23;
  reg  _T_84_isZero; // @[Reg.scala 11:16]
  reg [31:0] _RAND_24;
  reg  _T_84_sign; // @[Reg.scala 11:16]
  reg [31:0] _RAND_25;
  reg [12:0] _T_84_sExp; // @[Reg.scala 11:16]
  reg [31:0] _RAND_26;
  reg [55:0] _T_84_sig; // @[Reg.scala 11:16]
  reg [63:0] _RAND_27;
  reg [2:0] _T_93; // @[Reg.scala 11:16]
  reg [31:0] _RAND_28;
  reg  _T_102; // @[Reg.scala 11:16]
  reg [31:0] _RAND_29;
  reg  _T_109; // @[Valid.scala 48:22]
  reg [31:0] _RAND_30;
  reg  MulAddRecFNPipe_1_state; // @[Register tracking MulAddRecFNPipe_1 state]
  reg [31:0] _RAND_31;
  reg  MulAddRecFNPipe_1_cov [0:1]; // @[Coverage map for MulAddRecFNPipe_1]
  reg [31:0] _RAND_32;
  wire  MulAddRecFNPipe_1_cov_read_data; // @[Coverage map for MulAddRecFNPipe_1]
  wire  MulAddRecFNPipe_1_cov_read_addr; // @[Coverage map for MulAddRecFNPipe_1]
  wire  MulAddRecFNPipe_1_cov_write_data; // @[Coverage map for MulAddRecFNPipe_1]
  wire  MulAddRecFNPipe_1_cov_write_addr; // @[Coverage map for MulAddRecFNPipe_1]
  wire  MulAddRecFNPipe_1_cov_write_mask; // @[Coverage map for MulAddRecFNPipe_1]
  wire  MulAddRecFNPipe_1_cov_write_en; // @[Coverage map for MulAddRecFNPipe_1]
  reg [29:0] MulAddRecFNPipe_1_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_33;
  wire  valid_stage0_shl;
  wire  valid_stage0_pad;
  wire [29:0] mulAddRecFNToRaw_preMul_sum;
  wire [29:0] mulAddRecFNToRaw_postMul_sum;
  wire [29:0] roundRawFNToRecFN_sum;
  wire  mulAddRecFNToRaw_preMul_metaAssert_wire;
  wire  mulAddRecFNToRaw_postMul_metaAssert_wire;
  wire  roundRawFNToRecFN_metaAssert_wire;
  wire  MulAddRecFNPipe_1_or2;
  wire  MulAddRecFNPipe_1_or0;
  reg  MulAddRecFNPipe_1_metaAssert;
  reg [31:0] _RAND_34;
  MulAddRecFNToRaw_preMul_1 mulAddRecFNToRaw_preMul ( // @[FPU.scala 580:15]
    .io_op(mulAddRecFNToRaw_preMul_io_op),
    .io_a(mulAddRecFNToRaw_preMul_io_a),
    .io_b(mulAddRecFNToRaw_preMul_io_b),
    .io_c(mulAddRecFNToRaw_preMul_io_c),
    .io_mulAddA(mulAddRecFNToRaw_preMul_io_mulAddA),
    .io_mulAddB(mulAddRecFNToRaw_preMul_io_mulAddB),
    .io_mulAddC(mulAddRecFNToRaw_preMul_io_mulAddC),
    .io_toPostMul_isSigNaNAny(mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny),
    .io_toPostMul_isNaNAOrB(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB),
    .io_toPostMul_isInfA(mulAddRecFNToRaw_preMul_io_toPostMul_isInfA),
    .io_toPostMul_isZeroA(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA),
    .io_toPostMul_isInfB(mulAddRecFNToRaw_preMul_io_toPostMul_isInfB),
    .io_toPostMul_isZeroB(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB),
    .io_toPostMul_signProd(mulAddRecFNToRaw_preMul_io_toPostMul_signProd),
    .io_toPostMul_isNaNC(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC),
    .io_toPostMul_isInfC(mulAddRecFNToRaw_preMul_io_toPostMul_isInfC),
    .io_toPostMul_isZeroC(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC),
    .io_toPostMul_sExpSum(mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum),
    .io_toPostMul_doSubMags(mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags),
    .io_toPostMul_CIsDominant(mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant),
    .io_toPostMul_CDom_CAlignDist(mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist),
    .io_toPostMul_highAlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC),
    .io_toPostMul_bit0AlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC),
    .io_covSum(mulAddRecFNToRaw_preMul_io_covSum),
    .metaAssert(mulAddRecFNToRaw_preMul_metaAssert)
  );
  MulAddRecFNToRaw_postMul_1 mulAddRecFNToRaw_postMul ( // @[FPU.scala 582:15]
    .io_fromPreMul_isSigNaNAny(mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny),
    .io_fromPreMul_isNaNAOrB(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB),
    .io_fromPreMul_isInfA(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA),
    .io_fromPreMul_isZeroA(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA),
    .io_fromPreMul_isInfB(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB),
    .io_fromPreMul_isZeroB(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB),
    .io_fromPreMul_signProd(mulAddRecFNToRaw_postMul_io_fromPreMul_signProd),
    .io_fromPreMul_isNaNC(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC),
    .io_fromPreMul_isInfC(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC),
    .io_fromPreMul_isZeroC(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC),
    .io_fromPreMul_sExpSum(mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum),
    .io_fromPreMul_doSubMags(mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags),
    .io_fromPreMul_CIsDominant(mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant),
    .io_fromPreMul_CDom_CAlignDist(mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist),
    .io_fromPreMul_highAlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC),
    .io_fromPreMul_bit0AlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC),
    .io_mulAddResult(mulAddRecFNToRaw_postMul_io_mulAddResult),
    .io_roundingMode(mulAddRecFNToRaw_postMul_io_roundingMode),
    .io_invalidExc(mulAddRecFNToRaw_postMul_io_invalidExc),
    .io_rawOut_isNaN(mulAddRecFNToRaw_postMul_io_rawOut_isNaN),
    .io_rawOut_isInf(mulAddRecFNToRaw_postMul_io_rawOut_isInf),
    .io_rawOut_isZero(mulAddRecFNToRaw_postMul_io_rawOut_isZero),
    .io_rawOut_sign(mulAddRecFNToRaw_postMul_io_rawOut_sign),
    .io_rawOut_sExp(mulAddRecFNToRaw_postMul_io_rawOut_sExp),
    .io_rawOut_sig(mulAddRecFNToRaw_postMul_io_rawOut_sig),
    .io_covSum(mulAddRecFNToRaw_postMul_io_covSum),
    .metaAssert(mulAddRecFNToRaw_postMul_metaAssert)
  );
  RoundRawFNToRecFN_3 roundRawFNToRecFN ( // @[FPU.scala 608:35]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_infiniteExc(roundRawFNToRecFN_io_infiniteExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundRawFNToRecFN_io_detectTininess),
    .io_out(roundRawFNToRecFN_io_out),
    .io_exceptionFlags(roundRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundRawFNToRecFN_io_covSum),
    .metaAssert(roundRawFNToRecFN_metaAssert)
  );
  assign _T_14 = mulAddRecFNToRaw_preMul_io_mulAddA * mulAddRecFNToRaw_preMul_io_mulAddB; // @[FPU.scala 590:45]
  assign mulAddResult = _T_14 + mulAddRecFNToRaw_preMul_io_mulAddC; // @[FPU.scala 591:50]
  assign io_out = roundRawFNToRecFN_io_out; // @[FPU.scala 619:23]
  assign io_exceptionFlags = roundRawFNToRecFN_io_exceptionFlags; // @[FPU.scala 620:23]
  assign io_validout = _T_109; // @[FPU.scala 615:45]
  assign mulAddRecFNToRaw_preMul_io_op = io_op; // @[FPU.scala 584:35]
  assign mulAddRecFNToRaw_preMul_io_a = io_a; // @[FPU.scala 585:35]
  assign mulAddRecFNToRaw_preMul_io_b = io_b; // @[FPU.scala 586:35]
  assign mulAddRecFNToRaw_preMul_io_c = io_c; // @[FPU.scala 587:35]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny = _T_21_isSigNaNAny; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB = _T_21_isNaNAOrB; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA = _T_21_isInfA; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA = _T_21_isZeroA; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB = _T_21_isInfB; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB = _T_21_isZeroB; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_signProd = _T_21_signProd; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC = _T_21_isNaNC; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC = _T_21_isInfC; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC = _T_21_isZeroC; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum = _T_21_sExpSum; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags = _T_21_doSubMags; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant = _T_21_CIsDominant; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist = _T_21_CDom_CAlignDist; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC = _T_21_highAlignedSigC; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC = _T_21_bit0AlignedSigC; // @[FPU.scala 599:46]
  assign mulAddRecFNToRaw_postMul_io_mulAddResult = _T_30; // @[FPU.scala 600:46]
  assign mulAddRecFNToRaw_postMul_io_roundingMode = _T_39; // @[FPU.scala 601:46]
  assign roundRawFNToRecFN_io_invalidExc = _T_75; // @[FPU.scala 611:45]
  assign roundRawFNToRecFN_io_infiniteExc = 1'h0; // @[FPU.scala 617:38]
  assign roundRawFNToRecFN_io_in_isNaN = _T_84_isNaN; // @[FPU.scala 612:45]
  assign roundRawFNToRecFN_io_in_isInf = _T_84_isInf; // @[FPU.scala 612:45]
  assign roundRawFNToRecFN_io_in_isZero = _T_84_isZero; // @[FPU.scala 612:45]
  assign roundRawFNToRecFN_io_in_sign = _T_84_sign; // @[FPU.scala 612:45]
  assign roundRawFNToRecFN_io_in_sExp = _T_84_sExp; // @[FPU.scala 612:45]
  assign roundRawFNToRecFN_io_in_sig = _T_84_sig; // @[FPU.scala 612:45]
  assign roundRawFNToRecFN_io_roundingMode = _T_93; // @[FPU.scala 613:45]
  assign roundRawFNToRecFN_io_detectTininess = _T_102; // @[FPU.scala 614:45]
  assign MulAddRecFNPipe_1_cov_read_addr = MulAddRecFNPipe_1_state;
  assign MulAddRecFNPipe_1_cov_read_data = MulAddRecFNPipe_1_cov[MulAddRecFNPipe_1_cov_read_addr]; // @[Coverage map for MulAddRecFNPipe_1]
  assign MulAddRecFNPipe_1_cov_write_data = 1'h1;
  assign MulAddRecFNPipe_1_cov_write_addr = MulAddRecFNPipe_1_state;
  assign MulAddRecFNPipe_1_cov_write_mask = 1'h1;
  assign MulAddRecFNPipe_1_cov_write_en = 1'h1;
  assign valid_stage0_shl = valid_stage0;
  assign valid_stage0_pad = valid_stage0_shl;
  assign mulAddRecFNToRaw_preMul_sum = MulAddRecFNPipe_1_covSum + mulAddRecFNToRaw_preMul_io_covSum;
  assign mulAddRecFNToRaw_postMul_sum = mulAddRecFNToRaw_preMul_sum + mulAddRecFNToRaw_postMul_io_covSum;
  assign roundRawFNToRecFN_sum = mulAddRecFNToRaw_postMul_sum + roundRawFNToRecFN_io_covSum;
  assign io_covSum = roundRawFNToRecFN_sum;
  assign mulAddRecFNToRaw_preMul_metaAssert_wire = mulAddRecFNToRaw_preMul_metaAssert;
  assign mulAddRecFNToRaw_postMul_metaAssert_wire = mulAddRecFNToRaw_postMul_metaAssert;
  assign roundRawFNToRecFN_metaAssert_wire = roundRawFNToRecFN_metaAssert;
  assign MulAddRecFNPipe_1_or2 = mulAddRecFNToRaw_postMul_metaAssert_wire | roundRawFNToRecFN_metaAssert_wire;
  assign MulAddRecFNPipe_1_or0 = mulAddRecFNToRaw_preMul_metaAssert_wire | MulAddRecFNPipe_1_or2;
  assign metaAssert = MulAddRecFNPipe_1_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_21_isSigNaNAny = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_21_isNaNAOrB = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_21_isInfA = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_21_isZeroA = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_21_isInfB = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_21_isZeroB = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_21_signProd = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_21_isNaNC = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_21_isInfC = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_21_isZeroC = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_21_sExpSum = _RAND_10[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_21_doSubMags = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_21_CIsDominant = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_21_CDom_CAlignDist = _RAND_13[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {2{`RANDOM}};
  _T_21_highAlignedSigC = _RAND_14[54:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_21_bit0AlignedSigC = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {4{`RANDOM}};
  _T_30 = _RAND_16[106:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_39 = _RAND_17[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  roundingMode_stage0 = _RAND_18[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  detectTininess_stage0 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  valid_stage0 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_75 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_84_isNaN = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_84_isInf = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_84_isZero = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_84_sign = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_84_sExp = _RAND_26[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {2{`RANDOM}};
  _T_84_sig = _RAND_27[55:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_93 = _RAND_28[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_102 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_109 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  MulAddRecFNPipe_1_state = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    MulAddRecFNPipe_1_cov[initvar] = _RAND_32[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  MulAddRecFNPipe_1_covSum = _RAND_33[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  MulAddRecFNPipe_1_metaAssert = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      _T_21_isSigNaNAny <= 1'h0;
    end else if (io_validin) begin
      _T_21_isSigNaNAny <= mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny;
    end
    if (metaReset) begin
      _T_21_isNaNAOrB <= 1'h0;
    end else if (io_validin) begin
      _T_21_isNaNAOrB <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB;
    end
    if (metaReset) begin
      _T_21_isInfA <= 1'h0;
    end else if (io_validin) begin
      _T_21_isInfA <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfA;
    end
    if (metaReset) begin
      _T_21_isZeroA <= 1'h0;
    end else if (io_validin) begin
      _T_21_isZeroA <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA;
    end
    if (metaReset) begin
      _T_21_isInfB <= 1'h0;
    end else if (io_validin) begin
      _T_21_isInfB <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfB;
    end
    if (metaReset) begin
      _T_21_isZeroB <= 1'h0;
    end else if (io_validin) begin
      _T_21_isZeroB <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB;
    end
    if (metaReset) begin
      _T_21_signProd <= 1'h0;
    end else if (io_validin) begin
      _T_21_signProd <= mulAddRecFNToRaw_preMul_io_toPostMul_signProd;
    end
    if (metaReset) begin
      _T_21_isNaNC <= 1'h0;
    end else if (io_validin) begin
      _T_21_isNaNC <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC;
    end
    if (metaReset) begin
      _T_21_isInfC <= 1'h0;
    end else if (io_validin) begin
      _T_21_isInfC <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfC;
    end
    if (metaReset) begin
      _T_21_isZeroC <= 1'h0;
    end else if (io_validin) begin
      _T_21_isZeroC <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC;
    end
    if (metaReset) begin
      _T_21_sExpSum <= 13'h0;
    end else if (io_validin) begin
      _T_21_sExpSum <= mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum;
    end
    if (metaReset) begin
      _T_21_doSubMags <= 1'h0;
    end else if (io_validin) begin
      _T_21_doSubMags <= mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags;
    end
    if (metaReset) begin
      _T_21_CIsDominant <= 1'h0;
    end else if (io_validin) begin
      _T_21_CIsDominant <= mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant;
    end
    if (metaReset) begin
      _T_21_CDom_CAlignDist <= 6'h0;
    end else if (io_validin) begin
      _T_21_CDom_CAlignDist <= mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist;
    end
    if (metaReset) begin
      _T_21_highAlignedSigC <= 55'h0;
    end else if (io_validin) begin
      _T_21_highAlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC;
    end
    if (metaReset) begin
      _T_21_bit0AlignedSigC <= 1'h0;
    end else if (io_validin) begin
      _T_21_bit0AlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC;
    end
    if (metaReset) begin
      _T_30 <= 107'h0;
    end else if (io_validin) begin
      _T_30 <= mulAddResult;
    end
    if (metaReset) begin
      _T_39 <= 3'h0;
    end else if (io_validin) begin
      _T_39 <= io_roundingMode;
    end
    if (metaReset) begin
      roundingMode_stage0 <= 3'h0;
    end else if (io_validin) begin
      roundingMode_stage0 <= io_roundingMode;
    end
    if (metaReset) begin
      detectTininess_stage0 <= 1'h0;
    end else begin
      detectTininess_stage0 <= io_validin | detectTininess_stage0;
    end
    if (metaReset) begin
      valid_stage0 <= 1'h0;
    end else if (reset) begin
      valid_stage0 <= 1'h0;
    end else begin
      valid_stage0 <= io_validin;
    end
    if (metaReset) begin
      _T_75 <= 1'h0;
    end else if (valid_stage0) begin
      _T_75 <= mulAddRecFNToRaw_postMul_io_invalidExc;
    end
    if (metaReset) begin
      _T_84_isNaN <= 1'h0;
    end else if (valid_stage0) begin
      _T_84_isNaN <= mulAddRecFNToRaw_postMul_io_rawOut_isNaN;
    end
    if (metaReset) begin
      _T_84_isInf <= 1'h0;
    end else if (valid_stage0) begin
      _T_84_isInf <= mulAddRecFNToRaw_postMul_io_rawOut_isInf;
    end
    if (metaReset) begin
      _T_84_isZero <= 1'h0;
    end else if (valid_stage0) begin
      _T_84_isZero <= mulAddRecFNToRaw_postMul_io_rawOut_isZero;
    end
    if (metaReset) begin
      _T_84_sign <= 1'h0;
    end else if (valid_stage0) begin
      _T_84_sign <= mulAddRecFNToRaw_postMul_io_rawOut_sign;
    end
    if (metaReset) begin
      _T_84_sExp <= 13'h0;
    end else if (valid_stage0) begin
      _T_84_sExp <= mulAddRecFNToRaw_postMul_io_rawOut_sExp;
    end
    if (metaReset) begin
      _T_84_sig <= 56'h0;
    end else if (valid_stage0) begin
      _T_84_sig <= mulAddRecFNToRaw_postMul_io_rawOut_sig;
    end
    if (metaReset) begin
      _T_93 <= 3'h0;
    end else if (valid_stage0) begin
      _T_93 <= roundingMode_stage0;
    end
    if (metaReset) begin
      _T_102 <= 1'h0;
    end else if (valid_stage0) begin
      _T_102 <= detectTininess_stage0;
    end
    if (metaReset) begin
      _T_109 <= 1'h0;
    end else if (reset) begin
      _T_109 <= 1'h0;
    end else begin
      _T_109 <= valid_stage0;
    end
    MulAddRecFNPipe_1_state <= valid_stage0_pad;
    if (!(MulAddRecFNPipe_1_cov_read_data)) begin
      MulAddRecFNPipe_1_covSum <= MulAddRecFNPipe_1_covSum + 1'h1;
    end
    if (metaReset) begin
      MulAddRecFNPipe_1_metaAssert <= 1'h0;
    end else begin
      MulAddRecFNPipe_1_metaAssert <= MulAddRecFNPipe_1_metaAssert | MulAddRecFNPipe_1_or0;
    end
  end
  always @(posedge clock) begin
    if(MulAddRecFNPipe_1_cov_write_en & MulAddRecFNPipe_1_cov_write_mask) begin
      MulAddRecFNPipe_1_cov[MulAddRecFNPipe_1_cov_write_addr] <= MulAddRecFNPipe_1_cov_write_data; // @[Coverage map for MulAddRecFNPipe_1]
    end
  end
endmodule
module DivSqrtRecFNToRaw_small(
  input         clock,
  input         reset,
  output        io_inReady,
  input         io_inValid,
  input         io_sqrtOp,
  input  [32:0] io_a,
  input  [32:0] io_b,
  input  [2:0]  io_roundingMode,
  output        io_rawOutValid_div,
  output        io_rawOutValid_sqrt,
  output [2:0]  io_roundingModeOut,
  output        io_invalidExc,
  output        io_infiniteExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [9:0]  io_rawOut_sExp,
  output [26:0] io_rawOut_sig,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [4:0] cycleNum; // @[DivSqrtRecFN_small.scala 73:29]
  reg [31:0] _RAND_0;
  reg  sqrtOp_Z; // @[DivSqrtRecFN_small.scala 75:29]
  reg [31:0] _RAND_1;
  reg  majorExc_Z; // @[DivSqrtRecFN_small.scala 76:29]
  reg [31:0] _RAND_2;
  reg  isNaN_Z; // @[DivSqrtRecFN_small.scala 78:29]
  reg [31:0] _RAND_3;
  reg  isInf_Z; // @[DivSqrtRecFN_small.scala 79:29]
  reg [31:0] _RAND_4;
  reg  isZero_Z; // @[DivSqrtRecFN_small.scala 80:29]
  reg [31:0] _RAND_5;
  reg  sign_Z; // @[DivSqrtRecFN_small.scala 81:29]
  reg [31:0] _RAND_6;
  reg [9:0] sExp_Z; // @[DivSqrtRecFN_small.scala 82:29]
  reg [31:0] _RAND_7;
  reg [22:0] fractB_Z; // @[DivSqrtRecFN_small.scala 83:29]
  reg [31:0] _RAND_8;
  reg [2:0] roundingMode_Z; // @[DivSqrtRecFN_small.scala 84:29]
  reg [31:0] _RAND_9;
  reg [25:0] rem_Z; // @[DivSqrtRecFN_small.scala 90:29]
  reg [31:0] _RAND_10;
  reg  notZeroRem_Z; // @[DivSqrtRecFN_small.scala 91:29]
  reg [31:0] _RAND_11;
  reg [25:0] sigX_Z; // @[DivSqrtRecFN_small.scala 92:29]
  reg [31:0] _RAND_12;
  wire  rawA_S_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_33; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA_S_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawA_S_isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawA_S_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawA_S_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [24:0] rawA_S_sig; // @[Cat.scala 30:58]
  wire  rawB_S_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_50; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB_S_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawB_S_isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawB_S_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawB_S_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [24:0] rawB_S_sig; // @[Cat.scala 30:58]
  wire  _T_63; // @[DivSqrtRecFN_small.scala 101:24]
  wire  _T_64; // @[DivSqrtRecFN_small.scala 101:59]
  wire  notSigNaNIn_invalidExc_S_div; // @[DivSqrtRecFN_small.scala 101:42]
  wire  _T_67; // @[DivSqrtRecFN_small.scala 103:24]
  wire  notSigNaNIn_invalidExc_S_sqrt; // @[DivSqrtRecFN_small.scala 103:43]
  wire  _T_70; // @[common.scala 81:46]
  wire  _T_71; // @[DivSqrtRecFN_small.scala 106:38]
  wire  _T_77; // @[common.scala 81:46]
  wire  _T_78; // @[DivSqrtRecFN_small.scala 107:38]
  wire  _T_79; // @[DivSqrtRecFN_small.scala 107:66]
  wire  _T_82; // @[DivSqrtRecFN_small.scala 109:33]
  wire  _T_83; // @[DivSqrtRecFN_small.scala 109:51]
  wire  _T_84; // @[DivSqrtRecFN_small.scala 108:46]
  wire  _T_85; // @[DivSqrtRecFN_small.scala 113:26]
  wire  _T_86; // @[DivSqrtRecFN_small.scala 114:26]
  wire  _T_87; // @[DivSqrtRecFN_small.scala 114:42]
  wire  _T_88; // @[DivSqrtRecFN_small.scala 116:63]
  wire  _T_89; // @[DivSqrtRecFN_small.scala 117:64]
  wire  _T_91; // @[DivSqrtRecFN_small.scala 118:45]
  wire  sign_S; // @[DivSqrtRecFN_small.scala 118:30]
  wire  _T_92; // @[DivSqrtRecFN_small.scala 120:39]
  wire  specialCaseA_S; // @[DivSqrtRecFN_small.scala 120:55]
  wire  _T_93; // @[DivSqrtRecFN_small.scala 121:39]
  wire  specialCaseB_S; // @[DivSqrtRecFN_small.scala 121:55]
  wire  normalCase_S_div; // @[DivSqrtRecFN_small.scala 122:45]
  wire  normalCase_S_sqrt; // @[DivSqrtRecFN_small.scala 123:46]
  wire  normalCase_S; // @[DivSqrtRecFN_small.scala 124:27]
  wire [8:0] _T_102; // @[DivSqrtRecFN_small.scala 128:71]
  wire [9:0] _GEN_13; // @[DivSqrtRecFN_small.scala 127:21]
  wire [10:0] sExpQuot_S_div; // @[DivSqrtRecFN_small.scala 127:21]
  wire  _T_103; // @[DivSqrtRecFN_small.scala 131:50]
  wire [3:0] _T_105; // @[DivSqrtRecFN_small.scala 131:16]
  wire [9:0] sSatExpQuot_S_div; // @[DivSqrtRecFN_small.scala 136:11]
  wire  evenSqrt_S; // @[DivSqrtRecFN_small.scala 138:32]
  wire  oddSqrt_S; // @[DivSqrtRecFN_small.scala 139:32]
  wire  idle; // @[DivSqrtRecFN_small.scala 143:26]
  wire  inReady; // @[DivSqrtRecFN_small.scala 144:29]
  wire  entering; // @[DivSqrtRecFN_small.scala 145:28]
  wire  entering_normalCase; // @[DivSqrtRecFN_small.scala 146:40]
  wire  _T_111; // @[DivSqrtRecFN_small.scala 148:32]
  wire  skipCycle2; // @[DivSqrtRecFN_small.scala 148:45]
  wire  _T_114; // @[DivSqrtRecFN_small.scala 150:18]
  wire  _T_116; // @[DivSqrtRecFN_small.scala 152:26]
  wire [4:0] _T_119; // @[DivSqrtRecFN_small.scala 155:24]
  wire [4:0] _T_120; // @[DivSqrtRecFN_small.scala 154:20]
  wire [4:0] _T_121; // @[DivSqrtRecFN_small.scala 153:16]
  wire [4:0] _GEN_14; // @[DivSqrtRecFN_small.scala 152:62]
  wire [4:0] _T_122; // @[DivSqrtRecFN_small.scala 152:62]
  wire  _T_125; // @[DivSqrtRecFN_small.scala 160:24]
  wire [4:0] _T_128; // @[DivSqrtRecFN_small.scala 160:50]
  wire [4:0] _T_129; // @[DivSqrtRecFN_small.scala 160:16]
  wire [4:0] _T_130; // @[DivSqrtRecFN_small.scala 159:15]
  wire  _T_132; // @[DivSqrtRecFN_small.scala 161:24]
  wire [4:0] _GEN_15; // @[DivSqrtRecFN_small.scala 160:70]
  wire [4:0] _T_134; // @[DivSqrtRecFN_small.scala 160:70]
  wire [8:0] _T_135; // @[DivSqrtRecFN_small.scala 179:29]
  wire [9:0] _T_136; // @[DivSqrtRecFN_small.scala 179:34]
  wire  _T_139; // @[DivSqrtRecFN_small.scala 184:31]
  wire  _T_142; // @[DivSqrtRecFN_small.scala 191:21]
  wire [25:0] _T_143; // @[DivSqrtRecFN_small.scala 191:47]
  wire [25:0] _T_144; // @[DivSqrtRecFN_small.scala 191:12]
  wire  _T_145; // @[DivSqrtRecFN_small.scala 192:21]
  wire [1:0] _T_149; // @[DivSqrtRecFN_small.scala 193:56]
  wire [24:0] _T_151; // @[DivSqrtRecFN_small.scala 194:44]
  wire [26:0] _T_152; // @[Cat.scala 30:58]
  wire [26:0] _T_153; // @[DivSqrtRecFN_small.scala 192:12]
  wire [26:0] _GEN_16; // @[DivSqrtRecFN_small.scala 191:61]
  wire [26:0] _T_154; // @[DivSqrtRecFN_small.scala 191:61]
  wire [26:0] _T_156; // @[DivSqrtRecFN_small.scala 198:29]
  wire [26:0] _T_157; // @[DivSqrtRecFN_small.scala 198:12]
  wire [26:0] rem; // @[DivSqrtRecFN_small.scala 197:11]
  wire [31:0] _T_158; // @[DivSqrtRecFN_small.scala 199:27]
  wire [29:0] bitMask; // @[DivSqrtRecFN_small.scala 199:38]
  wire  _T_160; // @[DivSqrtRecFN_small.scala 201:21]
  wire [25:0] _T_161; // @[DivSqrtRecFN_small.scala 201:47]
  wire [25:0] _T_162; // @[DivSqrtRecFN_small.scala 201:12]
  wire  _T_163; // @[DivSqrtRecFN_small.scala 202:21]
  wire [24:0] _T_164; // @[DivSqrtRecFN_small.scala 202:12]
  wire [25:0] _GEN_17; // @[DivSqrtRecFN_small.scala 201:79]
  wire [25:0] _T_165; // @[DivSqrtRecFN_small.scala 201:79]
  wire [25:0] _T_167; // @[DivSqrtRecFN_small.scala 203:12]
  wire [25:0] _T_168; // @[DivSqrtRecFN_small.scala 202:79]
  wire  _T_171; // @[DivSqrtRecFN_small.scala 204:23]
  wire [23:0] _T_172; // @[Cat.scala 30:58]
  wire [24:0] _T_173; // @[DivSqrtRecFN_small.scala 204:63]
  wire [24:0] _T_174; // @[DivSqrtRecFN_small.scala 204:12]
  wire [25:0] _GEN_18; // @[DivSqrtRecFN_small.scala 203:79]
  wire [25:0] _T_175; // @[DivSqrtRecFN_small.scala 203:79]
  wire  _T_177; // @[DivSqrtRecFN_small.scala 205:23]
  wire [26:0] _T_178; // @[DivSqrtRecFN_small.scala 205:44]
  wire [29:0] _GEN_19; // @[DivSqrtRecFN_small.scala 205:48]
  wire [29:0] _T_179; // @[DivSqrtRecFN_small.scala 205:48]
  wire [29:0] _T_180; // @[DivSqrtRecFN_small.scala 205:12]
  wire [29:0] _GEN_20; // @[DivSqrtRecFN_small.scala 204:79]
  wire [29:0] trialTerm; // @[DivSqrtRecFN_small.scala 204:79]
  wire [27:0] _T_181; // @[DivSqrtRecFN_small.scala 206:24]
  wire [30:0] _T_182; // @[DivSqrtRecFN_small.scala 206:41]
  wire [30:0] _GEN_21; // @[DivSqrtRecFN_small.scala 206:29]
  wire [30:0] trialRem; // @[DivSqrtRecFN_small.scala 206:29]
  wire  newBit; // @[DivSqrtRecFN_small.scala 207:27]
  wire  _T_185; // @[DivSqrtRecFN_small.scala 209:44]
  wire  _T_186; // @[DivSqrtRecFN_small.scala 209:31]
  wire [30:0] _T_187; // @[DivSqrtRecFN_small.scala 210:39]
  wire [30:0] _T_188; // @[DivSqrtRecFN_small.scala 210:21]
  wire [30:0] _GEN_10; // @[DivSqrtRecFN_small.scala 209:56]
  wire  _T_190; // @[DivSqrtRecFN_small.scala 212:45]
  wire  _T_191; // @[DivSqrtRecFN_small.scala 212:31]
  wire  _T_192; // @[DivSqrtRecFN_small.scala 213:35]
  wire [25:0] _T_195; // @[DivSqrtRecFN_small.scala 215:47]
  wire [25:0] _T_196; // @[DivSqrtRecFN_small.scala 215:16]
  wire  _T_197; // @[DivSqrtRecFN_small.scala 216:25]
  wire [24:0] _T_198; // @[DivSqrtRecFN_small.scala 216:16]
  wire [25:0] _GEN_22; // @[DivSqrtRecFN_small.scala 215:77]
  wire [25:0] _T_199; // @[DivSqrtRecFN_small.scala 215:77]
  wire [23:0] _T_201; // @[DivSqrtRecFN_small.scala 217:47]
  wire [23:0] _T_202; // @[DivSqrtRecFN_small.scala 217:16]
  wire [25:0] _GEN_23; // @[DivSqrtRecFN_small.scala 216:77]
  wire [25:0] _T_203; // @[DivSqrtRecFN_small.scala 216:77]
  wire [29:0] _GEN_24; // @[DivSqrtRecFN_small.scala 218:48]
  wire [29:0] _T_205; // @[DivSqrtRecFN_small.scala 218:48]
  wire [29:0] _T_206; // @[DivSqrtRecFN_small.scala 218:16]
  wire [29:0] _GEN_25; // @[DivSqrtRecFN_small.scala 217:77]
  wire [29:0] _T_207; // @[DivSqrtRecFN_small.scala 217:77]
  wire [29:0] _GEN_12; // @[DivSqrtRecFN_small.scala 212:57]
  wire  rawOutValid; // @[DivSqrtRecFN_small.scala 223:33]
  wire [26:0] _GEN_26; // @[DivSqrtRecFN_small.scala 235:35]
  reg [5:0] DivSqrtRecFNToRaw_small_state; // @[Register tracking DivSqrtRecFNToRaw_small state]
  reg [31:0] _RAND_13;
  reg  DivSqrtRecFNToRaw_small_cov [0:63]; // @[Coverage map for DivSqrtRecFNToRaw_small]
  reg [31:0] _RAND_14;
  wire  DivSqrtRecFNToRaw_small_cov_read_data; // @[Coverage map for DivSqrtRecFNToRaw_small]
  wire [5:0] DivSqrtRecFNToRaw_small_cov_read_addr; // @[Coverage map for DivSqrtRecFNToRaw_small]
  wire  DivSqrtRecFNToRaw_small_cov_write_data; // @[Coverage map for DivSqrtRecFNToRaw_small]
  wire [5:0] DivSqrtRecFNToRaw_small_cov_write_addr; // @[Coverage map for DivSqrtRecFNToRaw_small]
  wire  DivSqrtRecFNToRaw_small_cov_write_mask; // @[Coverage map for DivSqrtRecFNToRaw_small]
  wire  DivSqrtRecFNToRaw_small_cov_write_en; // @[Coverage map for DivSqrtRecFNToRaw_small]
  reg [29:0] DivSqrtRecFNToRaw_small_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_15;
  wire  sqrtOp_Z_shl;
  wire [5:0] sqrtOp_Z_pad;
  wire [5:0] cycleNum_shl;
  wire [5:0] cycleNum_pad;
  wire [5:0] DivSqrtRecFNToRaw_small_xor0;
  assign rawA_S_isZero = io_a[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_33 = io_a[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawA_S_isNaN = _T_33 & io_a[29]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawA_S_isInf = _T_33 & ~io_a[29]; // @[rawFloatFromRecFN.scala 56:33]
  assign rawA_S_sign = io_a[32]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawA_S_sExp = {1'b0,$signed(io_a[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawA_S_sig = {1'h0,~rawA_S_isZero,io_a[22:0]}; // @[Cat.scala 30:58]
  assign rawB_S_isZero = io_b[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_50 = io_b[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawB_S_isNaN = _T_50 & io_b[29]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawB_S_isInf = _T_50 & ~io_b[29]; // @[rawFloatFromRecFN.scala 56:33]
  assign rawB_S_sign = io_b[32]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawB_S_sExp = {1'b0,$signed(io_b[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawB_S_sig = {1'h0,~rawB_S_isZero,io_b[22:0]}; // @[Cat.scala 30:58]
  assign _T_63 = rawA_S_isZero & rawB_S_isZero; // @[DivSqrtRecFN_small.scala 101:24]
  assign _T_64 = rawA_S_isInf & rawB_S_isInf; // @[DivSqrtRecFN_small.scala 101:59]
  assign notSigNaNIn_invalidExc_S_div = _T_63 | _T_64; // @[DivSqrtRecFN_small.scala 101:42]
  assign _T_67 = ~rawA_S_isNaN & ~rawA_S_isZero; // @[DivSqrtRecFN_small.scala 103:24]
  assign notSigNaNIn_invalidExc_S_sqrt = _T_67 & rawA_S_sign; // @[DivSqrtRecFN_small.scala 103:43]
  assign _T_70 = rawA_S_isNaN & ~rawA_S_sig[22]; // @[common.scala 81:46]
  assign _T_71 = _T_70 | notSigNaNIn_invalidExc_S_sqrt; // @[DivSqrtRecFN_small.scala 106:38]
  assign _T_77 = rawB_S_isNaN & ~rawB_S_sig[22]; // @[common.scala 81:46]
  assign _T_78 = _T_70 | _T_77; // @[DivSqrtRecFN_small.scala 107:38]
  assign _T_79 = _T_78 | notSigNaNIn_invalidExc_S_div; // @[DivSqrtRecFN_small.scala 107:66]
  assign _T_82 = ~rawA_S_isNaN & ~rawA_S_isInf; // @[DivSqrtRecFN_small.scala 109:33]
  assign _T_83 = _T_82 & rawB_S_isZero; // @[DivSqrtRecFN_small.scala 109:51]
  assign _T_84 = _T_79 | _T_83; // @[DivSqrtRecFN_small.scala 108:46]
  assign _T_85 = rawA_S_isNaN | notSigNaNIn_invalidExc_S_sqrt; // @[DivSqrtRecFN_small.scala 113:26]
  assign _T_86 = rawA_S_isNaN | rawB_S_isNaN; // @[DivSqrtRecFN_small.scala 114:26]
  assign _T_87 = _T_86 | notSigNaNIn_invalidExc_S_div; // @[DivSqrtRecFN_small.scala 114:42]
  assign _T_88 = rawA_S_isInf | rawB_S_isZero; // @[DivSqrtRecFN_small.scala 116:63]
  assign _T_89 = rawA_S_isZero | rawB_S_isInf; // @[DivSqrtRecFN_small.scala 117:64]
  assign _T_91 = ~io_sqrtOp & rawB_S_sign; // @[DivSqrtRecFN_small.scala 118:45]
  assign sign_S = rawA_S_sign ^ _T_91; // @[DivSqrtRecFN_small.scala 118:30]
  assign _T_92 = rawA_S_isNaN | rawA_S_isInf; // @[DivSqrtRecFN_small.scala 120:39]
  assign specialCaseA_S = _T_92 | rawA_S_isZero; // @[DivSqrtRecFN_small.scala 120:55]
  assign _T_93 = rawB_S_isNaN | rawB_S_isInf; // @[DivSqrtRecFN_small.scala 121:39]
  assign specialCaseB_S = _T_93 | rawB_S_isZero; // @[DivSqrtRecFN_small.scala 121:55]
  assign normalCase_S_div = ~specialCaseA_S & ~specialCaseB_S; // @[DivSqrtRecFN_small.scala 122:45]
  assign normalCase_S_sqrt = ~specialCaseA_S & ~rawA_S_sign; // @[DivSqrtRecFN_small.scala 123:46]
  assign normalCase_S = io_sqrtOp ? normalCase_S_sqrt : normalCase_S_div; // @[DivSqrtRecFN_small.scala 124:27]
  assign _T_102 = {rawB_S_sExp[8],~rawB_S_sExp[7:0]}; // @[DivSqrtRecFN_small.scala 128:71]
  assign _GEN_13 = {{1{_T_102[8]}},_T_102}; // @[DivSqrtRecFN_small.scala 127:21]
  assign sExpQuot_S_div = $signed(rawA_S_sExp) + $signed(_GEN_13); // @[DivSqrtRecFN_small.scala 127:21]
  assign _T_103 = 11'sh1c0 <= $signed(sExpQuot_S_div); // @[DivSqrtRecFN_small.scala 131:50]
  assign _T_105 = _T_103 ? 4'h6 : sExpQuot_S_div[9:6]; // @[DivSqrtRecFN_small.scala 131:16]
  assign sSatExpQuot_S_div = {_T_105,sExpQuot_S_div[5:0]}; // @[DivSqrtRecFN_small.scala 136:11]
  assign evenSqrt_S = io_sqrtOp & ~rawA_S_sExp[0]; // @[DivSqrtRecFN_small.scala 138:32]
  assign oddSqrt_S = io_sqrtOp & rawA_S_sExp[0]; // @[DivSqrtRecFN_small.scala 139:32]
  assign idle = cycleNum == 5'h0; // @[DivSqrtRecFN_small.scala 143:26]
  assign inReady = cycleNum <= 5'h1; // @[DivSqrtRecFN_small.scala 144:29]
  assign entering = inReady & io_inValid; // @[DivSqrtRecFN_small.scala 145:28]
  assign entering_normalCase = entering & normalCase_S; // @[DivSqrtRecFN_small.scala 146:40]
  assign _T_111 = cycleNum == 5'h3; // @[DivSqrtRecFN_small.scala 148:32]
  assign skipCycle2 = _T_111 & sigX_Z[25]; // @[DivSqrtRecFN_small.scala 148:45]
  assign _T_114 = ~idle | io_inValid; // @[DivSqrtRecFN_small.scala 150:18]
  assign _T_116 = entering & ~normalCase_S; // @[DivSqrtRecFN_small.scala 152:26]
  assign _T_119 = rawA_S_sExp[0] ? 5'h18 : 5'h19; // @[DivSqrtRecFN_small.scala 155:24]
  assign _T_120 = io_sqrtOp ? _T_119 : 5'h1a; // @[DivSqrtRecFN_small.scala 154:20]
  assign _T_121 = entering_normalCase ? _T_120 : 5'h0; // @[DivSqrtRecFN_small.scala 153:16]
  assign _GEN_14 = {{4'd0}, _T_116}; // @[DivSqrtRecFN_small.scala 152:62]
  assign _T_122 = _GEN_14 | _T_121; // @[DivSqrtRecFN_small.scala 152:62]
  assign _T_125 = ~idle & ~skipCycle2; // @[DivSqrtRecFN_small.scala 160:24]
  assign _T_128 = cycleNum - 5'h1; // @[DivSqrtRecFN_small.scala 160:50]
  assign _T_129 = _T_125 ? _T_128 : 5'h0; // @[DivSqrtRecFN_small.scala 160:16]
  assign _T_130 = _T_122 | _T_129; // @[DivSqrtRecFN_small.scala 159:15]
  assign _T_132 = ~idle & skipCycle2; // @[DivSqrtRecFN_small.scala 161:24]
  assign _GEN_15 = {{4'd0}, _T_132}; // @[DivSqrtRecFN_small.scala 160:70]
  assign _T_134 = _T_130 | _GEN_15; // @[DivSqrtRecFN_small.scala 160:70]
  assign _T_135 = rawA_S_sExp[9:1]; // @[DivSqrtRecFN_small.scala 179:29]
  assign _T_136 = $signed(_T_135) + 9'sh80; // @[DivSqrtRecFN_small.scala 179:34]
  assign _T_139 = entering_normalCase & ~io_sqrtOp; // @[DivSqrtRecFN_small.scala 184:31]
  assign _T_142 = inReady & ~oddSqrt_S; // @[DivSqrtRecFN_small.scala 191:21]
  assign _T_143 = {rawA_S_sig, 1'h0}; // @[DivSqrtRecFN_small.scala 191:47]
  assign _T_144 = _T_142 ? _T_143 : 26'h0; // @[DivSqrtRecFN_small.scala 191:12]
  assign _T_145 = inReady & oddSqrt_S; // @[DivSqrtRecFN_small.scala 192:21]
  assign _T_149 = rawA_S_sig[23:22] - 2'h1; // @[DivSqrtRecFN_small.scala 193:56]
  assign _T_151 = {rawA_S_sig[21:0], 3'h0}; // @[DivSqrtRecFN_small.scala 194:44]
  assign _T_152 = {_T_149,_T_151}; // @[Cat.scala 30:58]
  assign _T_153 = _T_145 ? _T_152 : 27'h0; // @[DivSqrtRecFN_small.scala 192:12]
  assign _GEN_16 = {{1'd0}, _T_144}; // @[DivSqrtRecFN_small.scala 191:61]
  assign _T_154 = _GEN_16 | _T_153; // @[DivSqrtRecFN_small.scala 191:61]
  assign _T_156 = {rem_Z, 1'h0}; // @[DivSqrtRecFN_small.scala 198:29]
  assign _T_157 = inReady ? 27'h0 : _T_156; // @[DivSqrtRecFN_small.scala 198:12]
  assign rem = _T_154 | _T_157; // @[DivSqrtRecFN_small.scala 197:11]
  assign _T_158 = 32'h1 << cycleNum; // @[DivSqrtRecFN_small.scala 199:27]
  assign bitMask = _T_158[31:2]; // @[DivSqrtRecFN_small.scala 199:38]
  assign _T_160 = inReady & ~io_sqrtOp; // @[DivSqrtRecFN_small.scala 201:21]
  assign _T_161 = {rawB_S_sig, 1'h0}; // @[DivSqrtRecFN_small.scala 201:47]
  assign _T_162 = _T_160 ? _T_161 : 26'h0; // @[DivSqrtRecFN_small.scala 201:12]
  assign _T_163 = inReady & evenSqrt_S; // @[DivSqrtRecFN_small.scala 202:21]
  assign _T_164 = _T_163 ? 25'h1000000 : 25'h0; // @[DivSqrtRecFN_small.scala 202:12]
  assign _GEN_17 = {{1'd0}, _T_164}; // @[DivSqrtRecFN_small.scala 201:79]
  assign _T_165 = _T_162 | _GEN_17; // @[DivSqrtRecFN_small.scala 201:79]
  assign _T_167 = _T_145 ? 26'h2800000 : 26'h0; // @[DivSqrtRecFN_small.scala 203:12]
  assign _T_168 = _T_165 | _T_167; // @[DivSqrtRecFN_small.scala 202:79]
  assign _T_171 = ~inReady & ~sqrtOp_Z; // @[DivSqrtRecFN_small.scala 204:23]
  assign _T_172 = {1'h1,fractB_Z}; // @[Cat.scala 30:58]
  assign _T_173 = {_T_172, 1'h0}; // @[DivSqrtRecFN_small.scala 204:63]
  assign _T_174 = _T_171 ? _T_173 : 25'h0; // @[DivSqrtRecFN_small.scala 204:12]
  assign _GEN_18 = {{1'd0}, _T_174}; // @[DivSqrtRecFN_small.scala 203:79]
  assign _T_175 = _T_168 | _GEN_18; // @[DivSqrtRecFN_small.scala 203:79]
  assign _T_177 = ~inReady & sqrtOp_Z; // @[DivSqrtRecFN_small.scala 205:23]
  assign _T_178 = {sigX_Z, 1'h0}; // @[DivSqrtRecFN_small.scala 205:44]
  assign _GEN_19 = {{3'd0}, _T_178}; // @[DivSqrtRecFN_small.scala 205:48]
  assign _T_179 = _GEN_19 | bitMask; // @[DivSqrtRecFN_small.scala 205:48]
  assign _T_180 = _T_177 ? _T_179 : 30'h0; // @[DivSqrtRecFN_small.scala 205:12]
  assign _GEN_20 = {{4'd0}, _T_175}; // @[DivSqrtRecFN_small.scala 204:79]
  assign trialTerm = _GEN_20 | _T_180; // @[DivSqrtRecFN_small.scala 204:79]
  assign _T_181 = {1'b0,$signed(rem)}; // @[DivSqrtRecFN_small.scala 206:24]
  assign _T_182 = {1'b0,$signed(trialTerm)}; // @[DivSqrtRecFN_small.scala 206:41]
  assign _GEN_21 = {{3{_T_181[27]}},_T_181}; // @[DivSqrtRecFN_small.scala 206:29]
  assign trialRem = $signed(_GEN_21) - $signed(_T_182); // @[DivSqrtRecFN_small.scala 206:29]
  assign newBit = 31'sh0 <= $signed(trialRem); // @[DivSqrtRecFN_small.scala 207:27]
  assign _T_185 = cycleNum > 5'h2; // @[DivSqrtRecFN_small.scala 209:44]
  assign _T_186 = entering_normalCase | _T_185; // @[DivSqrtRecFN_small.scala 209:31]
  assign _T_187 = $signed(_GEN_21) - $signed(_T_182); // @[DivSqrtRecFN_small.scala 210:39]
  assign _T_188 = newBit ? _T_187 : {{4'd0}, rem}; // @[DivSqrtRecFN_small.scala 210:21]
  assign _GEN_10 = _T_186 ? _T_188 : {{5'd0}, rem_Z}; // @[DivSqrtRecFN_small.scala 209:56]
  assign _T_190 = ~inReady & newBit; // @[DivSqrtRecFN_small.scala 212:45]
  assign _T_191 = entering_normalCase | _T_190; // @[DivSqrtRecFN_small.scala 212:31]
  assign _T_192 = $signed(trialRem) != 31'sh0; // @[DivSqrtRecFN_small.scala 213:35]
  assign _T_195 = {newBit, 25'h0}; // @[DivSqrtRecFN_small.scala 215:47]
  assign _T_196 = _T_160 ? _T_195 : 26'h0; // @[DivSqrtRecFN_small.scala 215:16]
  assign _T_197 = inReady & io_sqrtOp; // @[DivSqrtRecFN_small.scala 216:25]
  assign _T_198 = _T_197 ? 25'h1000000 : 25'h0; // @[DivSqrtRecFN_small.scala 216:16]
  assign _GEN_22 = {{1'd0}, _T_198}; // @[DivSqrtRecFN_small.scala 215:77]
  assign _T_199 = _T_196 | _GEN_22; // @[DivSqrtRecFN_small.scala 215:77]
  assign _T_201 = {newBit, 23'h0}; // @[DivSqrtRecFN_small.scala 217:47]
  assign _T_202 = _T_145 ? _T_201 : 24'h0; // @[DivSqrtRecFN_small.scala 217:16]
  assign _GEN_23 = {{2'd0}, _T_202}; // @[DivSqrtRecFN_small.scala 216:77]
  assign _T_203 = _T_199 | _GEN_23; // @[DivSqrtRecFN_small.scala 216:77]
  assign _GEN_24 = {{4'd0}, sigX_Z}; // @[DivSqrtRecFN_small.scala 218:48]
  assign _T_205 = _GEN_24 | bitMask; // @[DivSqrtRecFN_small.scala 218:48]
  assign _T_206 = inReady ? 30'h0 : _T_205; // @[DivSqrtRecFN_small.scala 218:16]
  assign _GEN_25 = {{4'd0}, _T_203}; // @[DivSqrtRecFN_small.scala 217:77]
  assign _T_207 = _GEN_25 | _T_206; // @[DivSqrtRecFN_small.scala 217:77]
  assign _GEN_12 = _T_191 ? _T_207 : {{4'd0}, sigX_Z}; // @[DivSqrtRecFN_small.scala 212:57]
  assign rawOutValid = cycleNum == 5'h1; // @[DivSqrtRecFN_small.scala 223:33]
  assign _GEN_26 = {{26'd0}, notZeroRem_Z}; // @[DivSqrtRecFN_small.scala 235:35]
  assign io_inReady = cycleNum <= 5'h1; // @[DivSqrtRecFN_small.scala 164:16]
  assign io_rawOutValid_div = rawOutValid & ~sqrtOp_Z; // @[DivSqrtRecFN_small.scala 225:25]
  assign io_rawOutValid_sqrt = rawOutValid & sqrtOp_Z; // @[DivSqrtRecFN_small.scala 226:25]
  assign io_roundingModeOut = roundingMode_Z; // @[DivSqrtRecFN_small.scala 227:25]
  assign io_invalidExc = majorExc_Z & isNaN_Z; // @[DivSqrtRecFN_small.scala 228:22]
  assign io_infiniteExc = majorExc_Z & ~isNaN_Z; // @[DivSqrtRecFN_small.scala 229:22]
  assign io_rawOut_isNaN = isNaN_Z; // @[DivSqrtRecFN_small.scala 230:22]
  assign io_rawOut_isInf = isInf_Z; // @[DivSqrtRecFN_small.scala 231:22]
  assign io_rawOut_isZero = isZero_Z; // @[DivSqrtRecFN_small.scala 232:22]
  assign io_rawOut_sign = sign_Z; // @[DivSqrtRecFN_small.scala 233:22]
  assign io_rawOut_sExp = sExp_Z; // @[DivSqrtRecFN_small.scala 234:22]
  assign io_rawOut_sig = _T_178 | _GEN_26; // @[DivSqrtRecFN_small.scala 235:22]
  assign DivSqrtRecFNToRaw_small_cov_read_addr = DivSqrtRecFNToRaw_small_state;
  assign DivSqrtRecFNToRaw_small_cov_read_data = DivSqrtRecFNToRaw_small_cov[DivSqrtRecFNToRaw_small_cov_read_addr]; // @[Coverage map for DivSqrtRecFNToRaw_small]
  assign DivSqrtRecFNToRaw_small_cov_write_data = 1'h1;
  assign DivSqrtRecFNToRaw_small_cov_write_addr = DivSqrtRecFNToRaw_small_state;
  assign DivSqrtRecFNToRaw_small_cov_write_mask = 1'h1;
  assign DivSqrtRecFNToRaw_small_cov_write_en = 1'h1;
  assign sqrtOp_Z_shl = sqrtOp_Z;
  assign sqrtOp_Z_pad = {5'h0,sqrtOp_Z_shl};
  assign cycleNum_shl = {cycleNum, 1'h0};
  assign cycleNum_pad = cycleNum_shl;
  assign DivSqrtRecFNToRaw_small_xor0 = sqrtOp_Z_pad ^ cycleNum_pad;
  assign io_covSum = DivSqrtRecFNToRaw_small_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleNum = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sqrtOp_Z = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  majorExc_Z = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  isNaN_Z = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  isInf_Z = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  isZero_Z = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sign_Z = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  sExp_Z = _RAND_7[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  fractB_Z = _RAND_8[22:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  roundingMode_Z = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  rem_Z = _RAND_10[25:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  notZeroRem_Z = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  sigX_Z = _RAND_12[25:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  DivSqrtRecFNToRaw_small_state = _RAND_13[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    DivSqrtRecFNToRaw_small_cov[initvar] = _RAND_14[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  DivSqrtRecFNToRaw_small_covSum = _RAND_15[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      cycleNum <= 5'h0;
    end else if (reset) begin
      cycleNum <= 5'h0;
    end else if (_T_114) begin
      cycleNum <= _T_134;
    end
    if (metaReset) begin
      sqrtOp_Z <= 1'h0;
    end else if (entering) begin
      sqrtOp_Z <= io_sqrtOp;
    end
    if (metaReset) begin
      majorExc_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        majorExc_Z <= _T_71;
      end else begin
        majorExc_Z <= _T_84;
      end
    end
    if (metaReset) begin
      isNaN_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        isNaN_Z <= _T_85;
      end else begin
        isNaN_Z <= _T_87;
      end
    end
    if (metaReset) begin
      isInf_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        isInf_Z <= rawA_S_isInf;
      end else begin
        isInf_Z <= _T_88;
      end
    end
    if (metaReset) begin
      isZero_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        isZero_Z <= rawA_S_isZero;
      end else begin
        isZero_Z <= _T_89;
      end
    end
    if (metaReset) begin
      sign_Z <= 1'h0;
    end else if (entering) begin
      sign_Z <= sign_S;
    end
    if (metaReset) begin
      sExp_Z <= 10'h0;
    end else if (entering_normalCase) begin
      if (io_sqrtOp) begin
        sExp_Z <= _T_136;
      end else begin
        sExp_Z <= sSatExpQuot_S_div;
      end
    end
    if (metaReset) begin
      fractB_Z <= 23'h0;
    end else if (_T_139) begin
      fractB_Z <= rawB_S_sig[22:0];
    end
    if (metaReset) begin
      roundingMode_Z <= 3'h0;
    end else if (entering_normalCase) begin
      roundingMode_Z <= io_roundingMode;
    end
    if (metaReset) begin
      rem_Z <= 26'h0;
    end else begin
      rem_Z <= _GEN_10[25:0];
    end
    if (metaReset) begin
      notZeroRem_Z <= 1'h0;
    end else if (_T_191) begin
      notZeroRem_Z <= _T_192;
    end
    if (metaReset) begin
      sigX_Z <= 26'h0;
    end else begin
      sigX_Z <= _GEN_12[25:0];
    end
    DivSqrtRecFNToRaw_small_state <= DivSqrtRecFNToRaw_small_xor0;
    if (!(DivSqrtRecFNToRaw_small_cov_read_data)) begin
      DivSqrtRecFNToRaw_small_covSum <= DivSqrtRecFNToRaw_small_covSum + 1'h1;
    end
  end
  always @(posedge clock) begin
    if(DivSqrtRecFNToRaw_small_cov_write_en & DivSqrtRecFNToRaw_small_cov_write_mask) begin
      DivSqrtRecFNToRaw_small_cov[DivSqrtRecFNToRaw_small_cov_write_addr] <= DivSqrtRecFNToRaw_small_cov_write_data; // @[Coverage map for DivSqrtRecFNToRaw_small]
    end
  end
endmodule
module RoundRawFNToRecFN_2(
  input         io_invalidExc,
  input         io_infiniteExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [9:0]  io_in_sExp,
  input  [26:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundAnyRawFNToRecFN_io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_infiniteExc; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [9:0] roundAnyRawFNToRecFN_io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [26:0] roundAnyRawFNToRecFN_io_in_sig; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [2:0] roundAnyRawFNToRecFN_io_roundingMode; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_detectTininess; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [32:0] roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [29:0] roundAnyRawFNToRecFN_io_covSum; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_metaAssert; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [29:0] RoundRawFNToRecFN_2_covSum;
  wire [29:0] roundAnyRawFNToRecFN_sum;
  wire  roundAnyRawFNToRecFN_metaAssert_wire;
  RoundAnyRawFNToRecFN_5 roundAnyRawFNToRecFN ( // @[RoundAnyRawFNToRecFN.scala 307:15]
    .io_invalidExc(roundAnyRawFNToRecFN_io_invalidExc),
    .io_infiniteExc(roundAnyRawFNToRecFN_io_infiniteExc),
    .io_in_isNaN(roundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundAnyRawFNToRecFN_io_detectTininess),
    .io_out(roundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundAnyRawFNToRecFN_io_covSum),
    .metaAssert(roundAnyRawFNToRecFN_metaAssert)
  );
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 315:23]
  assign io_exceptionFlags = roundAnyRawFNToRecFN_io_exceptionFlags; // @[RoundAnyRawFNToRecFN.scala 316:23]
  assign roundAnyRawFNToRecFN_io_invalidExc = io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 310:44]
  assign roundAnyRawFNToRecFN_io_infiniteExc = io_infiniteExc; // @[RoundAnyRawFNToRecFN.scala 311:44]
  assign roundAnyRawFNToRecFN_io_in_isNaN = io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isInf = io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isZero = io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_in_sign; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sig = io_in_sig; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[RoundAnyRawFNToRecFN.scala 313:44]
  assign roundAnyRawFNToRecFN_io_detectTininess = io_detectTininess; // @[RoundAnyRawFNToRecFN.scala 314:44]
  assign RoundRawFNToRecFN_2_covSum = 30'h0;
  assign roundAnyRawFNToRecFN_sum = RoundRawFNToRecFN_2_covSum + roundAnyRawFNToRecFN_io_covSum;
  assign io_covSum = roundAnyRawFNToRecFN_sum;
  assign roundAnyRawFNToRecFN_metaAssert_wire = roundAnyRawFNToRecFN_metaAssert;
  assign metaAssert = roundAnyRawFNToRecFN_metaAssert_wire;
endmodule
module DivSqrtRecFNToRaw_small_1(
  input         clock,
  input         reset,
  output        io_inReady,
  input         io_inValid,
  input         io_sqrtOp,
  input  [64:0] io_a,
  input  [64:0] io_b,
  input  [2:0]  io_roundingMode,
  output        io_rawOutValid_div,
  output        io_rawOutValid_sqrt,
  output [2:0]  io_roundingModeOut,
  output        io_invalidExc,
  output        io_infiniteExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [12:0] io_rawOut_sExp,
  output [55:0] io_rawOut_sig,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [5:0] cycleNum; // @[DivSqrtRecFN_small.scala 73:29]
  reg [31:0] _RAND_0;
  reg  sqrtOp_Z; // @[DivSqrtRecFN_small.scala 75:29]
  reg [31:0] _RAND_1;
  reg  majorExc_Z; // @[DivSqrtRecFN_small.scala 76:29]
  reg [31:0] _RAND_2;
  reg  isNaN_Z; // @[DivSqrtRecFN_small.scala 78:29]
  reg [31:0] _RAND_3;
  reg  isInf_Z; // @[DivSqrtRecFN_small.scala 79:29]
  reg [31:0] _RAND_4;
  reg  isZero_Z; // @[DivSqrtRecFN_small.scala 80:29]
  reg [31:0] _RAND_5;
  reg  sign_Z; // @[DivSqrtRecFN_small.scala 81:29]
  reg [31:0] _RAND_6;
  reg [12:0] sExp_Z; // @[DivSqrtRecFN_small.scala 82:29]
  reg [31:0] _RAND_7;
  reg [51:0] fractB_Z; // @[DivSqrtRecFN_small.scala 83:29]
  reg [63:0] _RAND_8;
  reg [2:0] roundingMode_Z; // @[DivSqrtRecFN_small.scala 84:29]
  reg [31:0] _RAND_9;
  reg [54:0] rem_Z; // @[DivSqrtRecFN_small.scala 90:29]
  reg [63:0] _RAND_10;
  reg  notZeroRem_Z; // @[DivSqrtRecFN_small.scala 91:29]
  reg [31:0] _RAND_11;
  reg [54:0] sigX_Z; // @[DivSqrtRecFN_small.scala 92:29]
  reg [63:0] _RAND_12;
  wire  rawA_S_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_33; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA_S_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawA_S_isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawA_S_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawA_S_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] rawA_S_sig; // @[Cat.scala 30:58]
  wire  rawB_S_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_50; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB_S_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawB_S_isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawB_S_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawB_S_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] rawB_S_sig; // @[Cat.scala 30:58]
  wire  _T_63; // @[DivSqrtRecFN_small.scala 101:24]
  wire  _T_64; // @[DivSqrtRecFN_small.scala 101:59]
  wire  notSigNaNIn_invalidExc_S_div; // @[DivSqrtRecFN_small.scala 101:42]
  wire  _T_67; // @[DivSqrtRecFN_small.scala 103:24]
  wire  notSigNaNIn_invalidExc_S_sqrt; // @[DivSqrtRecFN_small.scala 103:43]
  wire  _T_70; // @[common.scala 81:46]
  wire  _T_71; // @[DivSqrtRecFN_small.scala 106:38]
  wire  _T_77; // @[common.scala 81:46]
  wire  _T_78; // @[DivSqrtRecFN_small.scala 107:38]
  wire  _T_79; // @[DivSqrtRecFN_small.scala 107:66]
  wire  _T_82; // @[DivSqrtRecFN_small.scala 109:33]
  wire  _T_83; // @[DivSqrtRecFN_small.scala 109:51]
  wire  _T_84; // @[DivSqrtRecFN_small.scala 108:46]
  wire  _T_85; // @[DivSqrtRecFN_small.scala 113:26]
  wire  _T_86; // @[DivSqrtRecFN_small.scala 114:26]
  wire  _T_87; // @[DivSqrtRecFN_small.scala 114:42]
  wire  _T_88; // @[DivSqrtRecFN_small.scala 116:63]
  wire  _T_89; // @[DivSqrtRecFN_small.scala 117:64]
  wire  _T_91; // @[DivSqrtRecFN_small.scala 118:45]
  wire  sign_S; // @[DivSqrtRecFN_small.scala 118:30]
  wire  _T_92; // @[DivSqrtRecFN_small.scala 120:39]
  wire  specialCaseA_S; // @[DivSqrtRecFN_small.scala 120:55]
  wire  _T_93; // @[DivSqrtRecFN_small.scala 121:39]
  wire  specialCaseB_S; // @[DivSqrtRecFN_small.scala 121:55]
  wire  normalCase_S_div; // @[DivSqrtRecFN_small.scala 122:45]
  wire  normalCase_S_sqrt; // @[DivSqrtRecFN_small.scala 123:46]
  wire  normalCase_S; // @[DivSqrtRecFN_small.scala 124:27]
  wire [11:0] _T_102; // @[DivSqrtRecFN_small.scala 128:71]
  wire [12:0] _GEN_13; // @[DivSqrtRecFN_small.scala 127:21]
  wire [13:0] sExpQuot_S_div; // @[DivSqrtRecFN_small.scala 127:21]
  wire  _T_103; // @[DivSqrtRecFN_small.scala 131:50]
  wire [3:0] _T_105; // @[DivSqrtRecFN_small.scala 131:16]
  wire [12:0] sSatExpQuot_S_div; // @[DivSqrtRecFN_small.scala 136:11]
  wire  evenSqrt_S; // @[DivSqrtRecFN_small.scala 138:32]
  wire  oddSqrt_S; // @[DivSqrtRecFN_small.scala 139:32]
  wire  idle; // @[DivSqrtRecFN_small.scala 143:26]
  wire  inReady; // @[DivSqrtRecFN_small.scala 144:29]
  wire  entering; // @[DivSqrtRecFN_small.scala 145:28]
  wire  entering_normalCase; // @[DivSqrtRecFN_small.scala 146:40]
  wire  _T_111; // @[DivSqrtRecFN_small.scala 148:32]
  wire  skipCycle2; // @[DivSqrtRecFN_small.scala 148:45]
  wire  _T_114; // @[DivSqrtRecFN_small.scala 150:18]
  wire  _T_116; // @[DivSqrtRecFN_small.scala 152:26]
  wire [5:0] _T_119; // @[DivSqrtRecFN_small.scala 155:24]
  wire [5:0] _T_120; // @[DivSqrtRecFN_small.scala 154:20]
  wire [5:0] _T_121; // @[DivSqrtRecFN_small.scala 153:16]
  wire [5:0] _GEN_14; // @[DivSqrtRecFN_small.scala 152:62]
  wire [5:0] _T_122; // @[DivSqrtRecFN_small.scala 152:62]
  wire  _T_125; // @[DivSqrtRecFN_small.scala 160:24]
  wire [5:0] _T_128; // @[DivSqrtRecFN_small.scala 160:50]
  wire [5:0] _T_129; // @[DivSqrtRecFN_small.scala 160:16]
  wire [5:0] _T_130; // @[DivSqrtRecFN_small.scala 159:15]
  wire  _T_132; // @[DivSqrtRecFN_small.scala 161:24]
  wire [5:0] _GEN_15; // @[DivSqrtRecFN_small.scala 160:70]
  wire [5:0] _T_134; // @[DivSqrtRecFN_small.scala 160:70]
  wire [11:0] _T_135; // @[DivSqrtRecFN_small.scala 179:29]
  wire [12:0] _T_136; // @[DivSqrtRecFN_small.scala 179:34]
  wire  _T_139; // @[DivSqrtRecFN_small.scala 184:31]
  wire  _T_142; // @[DivSqrtRecFN_small.scala 191:21]
  wire [54:0] _T_143; // @[DivSqrtRecFN_small.scala 191:47]
  wire [54:0] _T_144; // @[DivSqrtRecFN_small.scala 191:12]
  wire  _T_145; // @[DivSqrtRecFN_small.scala 192:21]
  wire [1:0] _T_149; // @[DivSqrtRecFN_small.scala 193:56]
  wire [53:0] _T_151; // @[DivSqrtRecFN_small.scala 194:44]
  wire [55:0] _T_152; // @[Cat.scala 30:58]
  wire [55:0] _T_153; // @[DivSqrtRecFN_small.scala 192:12]
  wire [55:0] _GEN_16; // @[DivSqrtRecFN_small.scala 191:61]
  wire [55:0] _T_154; // @[DivSqrtRecFN_small.scala 191:61]
  wire [55:0] _T_156; // @[DivSqrtRecFN_small.scala 198:29]
  wire [55:0] _T_157; // @[DivSqrtRecFN_small.scala 198:12]
  wire [55:0] rem; // @[DivSqrtRecFN_small.scala 197:11]
  wire [63:0] _T_158; // @[DivSqrtRecFN_small.scala 199:27]
  wire [61:0] bitMask; // @[DivSqrtRecFN_small.scala 199:38]
  wire  _T_160; // @[DivSqrtRecFN_small.scala 201:21]
  wire [54:0] _T_161; // @[DivSqrtRecFN_small.scala 201:47]
  wire [54:0] _T_162; // @[DivSqrtRecFN_small.scala 201:12]
  wire  _T_163; // @[DivSqrtRecFN_small.scala 202:21]
  wire [53:0] _T_164; // @[DivSqrtRecFN_small.scala 202:12]
  wire [54:0] _GEN_17; // @[DivSqrtRecFN_small.scala 201:79]
  wire [54:0] _T_165; // @[DivSqrtRecFN_small.scala 201:79]
  wire [54:0] _T_167; // @[DivSqrtRecFN_small.scala 203:12]
  wire [54:0] _T_168; // @[DivSqrtRecFN_small.scala 202:79]
  wire  _T_171; // @[DivSqrtRecFN_small.scala 204:23]
  wire [52:0] _T_172; // @[Cat.scala 30:58]
  wire [53:0] _T_173; // @[DivSqrtRecFN_small.scala 204:63]
  wire [53:0] _T_174; // @[DivSqrtRecFN_small.scala 204:12]
  wire [54:0] _GEN_18; // @[DivSqrtRecFN_small.scala 203:79]
  wire [54:0] _T_175; // @[DivSqrtRecFN_small.scala 203:79]
  wire  _T_177; // @[DivSqrtRecFN_small.scala 205:23]
  wire [55:0] _T_178; // @[DivSqrtRecFN_small.scala 205:44]
  wire [61:0] _GEN_19; // @[DivSqrtRecFN_small.scala 205:48]
  wire [61:0] _T_179; // @[DivSqrtRecFN_small.scala 205:48]
  wire [61:0] _T_180; // @[DivSqrtRecFN_small.scala 205:12]
  wire [61:0] _GEN_20; // @[DivSqrtRecFN_small.scala 204:79]
  wire [61:0] trialTerm; // @[DivSqrtRecFN_small.scala 204:79]
  wire [56:0] _T_181; // @[DivSqrtRecFN_small.scala 206:24]
  wire [62:0] _T_182; // @[DivSqrtRecFN_small.scala 206:41]
  wire [62:0] _GEN_21; // @[DivSqrtRecFN_small.scala 206:29]
  wire [62:0] trialRem; // @[DivSqrtRecFN_small.scala 206:29]
  wire  newBit; // @[DivSqrtRecFN_small.scala 207:27]
  wire  _T_185; // @[DivSqrtRecFN_small.scala 209:44]
  wire  _T_186; // @[DivSqrtRecFN_small.scala 209:31]
  wire [62:0] _T_187; // @[DivSqrtRecFN_small.scala 210:39]
  wire [62:0] _T_188; // @[DivSqrtRecFN_small.scala 210:21]
  wire [62:0] _GEN_10; // @[DivSqrtRecFN_small.scala 209:56]
  wire  _T_190; // @[DivSqrtRecFN_small.scala 212:45]
  wire  _T_191; // @[DivSqrtRecFN_small.scala 212:31]
  wire  _T_192; // @[DivSqrtRecFN_small.scala 213:35]
  wire [54:0] _T_195; // @[DivSqrtRecFN_small.scala 215:47]
  wire [54:0] _T_196; // @[DivSqrtRecFN_small.scala 215:16]
  wire  _T_197; // @[DivSqrtRecFN_small.scala 216:25]
  wire [53:0] _T_198; // @[DivSqrtRecFN_small.scala 216:16]
  wire [54:0] _GEN_22; // @[DivSqrtRecFN_small.scala 215:77]
  wire [54:0] _T_199; // @[DivSqrtRecFN_small.scala 215:77]
  wire [52:0] _T_201; // @[DivSqrtRecFN_small.scala 217:47]
  wire [52:0] _T_202; // @[DivSqrtRecFN_small.scala 217:16]
  wire [54:0] _GEN_23; // @[DivSqrtRecFN_small.scala 216:77]
  wire [54:0] _T_203; // @[DivSqrtRecFN_small.scala 216:77]
  wire [61:0] _GEN_24; // @[DivSqrtRecFN_small.scala 218:48]
  wire [61:0] _T_205; // @[DivSqrtRecFN_small.scala 218:48]
  wire [61:0] _T_206; // @[DivSqrtRecFN_small.scala 218:16]
  wire [61:0] _GEN_25; // @[DivSqrtRecFN_small.scala 217:77]
  wire [61:0] _T_207; // @[DivSqrtRecFN_small.scala 217:77]
  wire [61:0] _GEN_12; // @[DivSqrtRecFN_small.scala 212:57]
  wire  rawOutValid; // @[DivSqrtRecFN_small.scala 223:33]
  wire [55:0] _GEN_26; // @[DivSqrtRecFN_small.scala 235:35]
  reg [6:0] DivSqrtRecFNToRaw_small_1_state; // @[Register tracking DivSqrtRecFNToRaw_small_1 state]
  reg [31:0] _RAND_13;
  reg  DivSqrtRecFNToRaw_small_1_cov [0:127]; // @[Coverage map for DivSqrtRecFNToRaw_small_1]
  reg [31:0] _RAND_14;
  wire  DivSqrtRecFNToRaw_small_1_cov_read_data; // @[Coverage map for DivSqrtRecFNToRaw_small_1]
  wire [6:0] DivSqrtRecFNToRaw_small_1_cov_read_addr; // @[Coverage map for DivSqrtRecFNToRaw_small_1]
  wire  DivSqrtRecFNToRaw_small_1_cov_write_data; // @[Coverage map for DivSqrtRecFNToRaw_small_1]
  wire [6:0] DivSqrtRecFNToRaw_small_1_cov_write_addr; // @[Coverage map for DivSqrtRecFNToRaw_small_1]
  wire  DivSqrtRecFNToRaw_small_1_cov_write_mask; // @[Coverage map for DivSqrtRecFNToRaw_small_1]
  wire  DivSqrtRecFNToRaw_small_1_cov_write_en; // @[Coverage map for DivSqrtRecFNToRaw_small_1]
  reg [29:0] DivSqrtRecFNToRaw_small_1_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_15;
  wire  sqrtOp_Z_shl;
  wire [6:0] sqrtOp_Z_pad;
  wire [6:0] cycleNum_shl;
  wire [6:0] cycleNum_pad;
  wire [6:0] DivSqrtRecFNToRaw_small_1_xor0;
  assign rawA_S_isZero = io_a[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_33 = io_a[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawA_S_isNaN = _T_33 & io_a[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawA_S_isInf = _T_33 & ~io_a[61]; // @[rawFloatFromRecFN.scala 56:33]
  assign rawA_S_sign = io_a[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawA_S_sExp = {1'b0,$signed(io_a[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawA_S_sig = {1'h0,~rawA_S_isZero,io_a[51:0]}; // @[Cat.scala 30:58]
  assign rawB_S_isZero = io_b[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_50 = io_b[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawB_S_isNaN = _T_50 & io_b[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawB_S_isInf = _T_50 & ~io_b[61]; // @[rawFloatFromRecFN.scala 56:33]
  assign rawB_S_sign = io_b[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawB_S_sExp = {1'b0,$signed(io_b[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawB_S_sig = {1'h0,~rawB_S_isZero,io_b[51:0]}; // @[Cat.scala 30:58]
  assign _T_63 = rawA_S_isZero & rawB_S_isZero; // @[DivSqrtRecFN_small.scala 101:24]
  assign _T_64 = rawA_S_isInf & rawB_S_isInf; // @[DivSqrtRecFN_small.scala 101:59]
  assign notSigNaNIn_invalidExc_S_div = _T_63 | _T_64; // @[DivSqrtRecFN_small.scala 101:42]
  assign _T_67 = ~rawA_S_isNaN & ~rawA_S_isZero; // @[DivSqrtRecFN_small.scala 103:24]
  assign notSigNaNIn_invalidExc_S_sqrt = _T_67 & rawA_S_sign; // @[DivSqrtRecFN_small.scala 103:43]
  assign _T_70 = rawA_S_isNaN & ~rawA_S_sig[51]; // @[common.scala 81:46]
  assign _T_71 = _T_70 | notSigNaNIn_invalidExc_S_sqrt; // @[DivSqrtRecFN_small.scala 106:38]
  assign _T_77 = rawB_S_isNaN & ~rawB_S_sig[51]; // @[common.scala 81:46]
  assign _T_78 = _T_70 | _T_77; // @[DivSqrtRecFN_small.scala 107:38]
  assign _T_79 = _T_78 | notSigNaNIn_invalidExc_S_div; // @[DivSqrtRecFN_small.scala 107:66]
  assign _T_82 = ~rawA_S_isNaN & ~rawA_S_isInf; // @[DivSqrtRecFN_small.scala 109:33]
  assign _T_83 = _T_82 & rawB_S_isZero; // @[DivSqrtRecFN_small.scala 109:51]
  assign _T_84 = _T_79 | _T_83; // @[DivSqrtRecFN_small.scala 108:46]
  assign _T_85 = rawA_S_isNaN | notSigNaNIn_invalidExc_S_sqrt; // @[DivSqrtRecFN_small.scala 113:26]
  assign _T_86 = rawA_S_isNaN | rawB_S_isNaN; // @[DivSqrtRecFN_small.scala 114:26]
  assign _T_87 = _T_86 | notSigNaNIn_invalidExc_S_div; // @[DivSqrtRecFN_small.scala 114:42]
  assign _T_88 = rawA_S_isInf | rawB_S_isZero; // @[DivSqrtRecFN_small.scala 116:63]
  assign _T_89 = rawA_S_isZero | rawB_S_isInf; // @[DivSqrtRecFN_small.scala 117:64]
  assign _T_91 = ~io_sqrtOp & rawB_S_sign; // @[DivSqrtRecFN_small.scala 118:45]
  assign sign_S = rawA_S_sign ^ _T_91; // @[DivSqrtRecFN_small.scala 118:30]
  assign _T_92 = rawA_S_isNaN | rawA_S_isInf; // @[DivSqrtRecFN_small.scala 120:39]
  assign specialCaseA_S = _T_92 | rawA_S_isZero; // @[DivSqrtRecFN_small.scala 120:55]
  assign _T_93 = rawB_S_isNaN | rawB_S_isInf; // @[DivSqrtRecFN_small.scala 121:39]
  assign specialCaseB_S = _T_93 | rawB_S_isZero; // @[DivSqrtRecFN_small.scala 121:55]
  assign normalCase_S_div = ~specialCaseA_S & ~specialCaseB_S; // @[DivSqrtRecFN_small.scala 122:45]
  assign normalCase_S_sqrt = ~specialCaseA_S & ~rawA_S_sign; // @[DivSqrtRecFN_small.scala 123:46]
  assign normalCase_S = io_sqrtOp ? normalCase_S_sqrt : normalCase_S_div; // @[DivSqrtRecFN_small.scala 124:27]
  assign _T_102 = {rawB_S_sExp[11],~rawB_S_sExp[10:0]}; // @[DivSqrtRecFN_small.scala 128:71]
  assign _GEN_13 = {{1{_T_102[11]}},_T_102}; // @[DivSqrtRecFN_small.scala 127:21]
  assign sExpQuot_S_div = $signed(rawA_S_sExp) + $signed(_GEN_13); // @[DivSqrtRecFN_small.scala 127:21]
  assign _T_103 = 14'she00 <= $signed(sExpQuot_S_div); // @[DivSqrtRecFN_small.scala 131:50]
  assign _T_105 = _T_103 ? 4'h6 : sExpQuot_S_div[12:9]; // @[DivSqrtRecFN_small.scala 131:16]
  assign sSatExpQuot_S_div = {_T_105,sExpQuot_S_div[8:0]}; // @[DivSqrtRecFN_small.scala 136:11]
  assign evenSqrt_S = io_sqrtOp & ~rawA_S_sExp[0]; // @[DivSqrtRecFN_small.scala 138:32]
  assign oddSqrt_S = io_sqrtOp & rawA_S_sExp[0]; // @[DivSqrtRecFN_small.scala 139:32]
  assign idle = cycleNum == 6'h0; // @[DivSqrtRecFN_small.scala 143:26]
  assign inReady = cycleNum <= 6'h1; // @[DivSqrtRecFN_small.scala 144:29]
  assign entering = inReady & io_inValid; // @[DivSqrtRecFN_small.scala 145:28]
  assign entering_normalCase = entering & normalCase_S; // @[DivSqrtRecFN_small.scala 146:40]
  assign _T_111 = cycleNum == 6'h3; // @[DivSqrtRecFN_small.scala 148:32]
  assign skipCycle2 = _T_111 & sigX_Z[54]; // @[DivSqrtRecFN_small.scala 148:45]
  assign _T_114 = ~idle | io_inValid; // @[DivSqrtRecFN_small.scala 150:18]
  assign _T_116 = entering & ~normalCase_S; // @[DivSqrtRecFN_small.scala 152:26]
  assign _T_119 = rawA_S_sExp[0] ? 6'h35 : 6'h36; // @[DivSqrtRecFN_small.scala 155:24]
  assign _T_120 = io_sqrtOp ? _T_119 : 6'h37; // @[DivSqrtRecFN_small.scala 154:20]
  assign _T_121 = entering_normalCase ? _T_120 : 6'h0; // @[DivSqrtRecFN_small.scala 153:16]
  assign _GEN_14 = {{5'd0}, _T_116}; // @[DivSqrtRecFN_small.scala 152:62]
  assign _T_122 = _GEN_14 | _T_121; // @[DivSqrtRecFN_small.scala 152:62]
  assign _T_125 = ~idle & ~skipCycle2; // @[DivSqrtRecFN_small.scala 160:24]
  assign _T_128 = cycleNum - 6'h1; // @[DivSqrtRecFN_small.scala 160:50]
  assign _T_129 = _T_125 ? _T_128 : 6'h0; // @[DivSqrtRecFN_small.scala 160:16]
  assign _T_130 = _T_122 | _T_129; // @[DivSqrtRecFN_small.scala 159:15]
  assign _T_132 = ~idle & skipCycle2; // @[DivSqrtRecFN_small.scala 161:24]
  assign _GEN_15 = {{5'd0}, _T_132}; // @[DivSqrtRecFN_small.scala 160:70]
  assign _T_134 = _T_130 | _GEN_15; // @[DivSqrtRecFN_small.scala 160:70]
  assign _T_135 = rawA_S_sExp[12:1]; // @[DivSqrtRecFN_small.scala 179:29]
  assign _T_136 = $signed(_T_135) + 12'sh400; // @[DivSqrtRecFN_small.scala 179:34]
  assign _T_139 = entering_normalCase & ~io_sqrtOp; // @[DivSqrtRecFN_small.scala 184:31]
  assign _T_142 = inReady & ~oddSqrt_S; // @[DivSqrtRecFN_small.scala 191:21]
  assign _T_143 = {rawA_S_sig, 1'h0}; // @[DivSqrtRecFN_small.scala 191:47]
  assign _T_144 = _T_142 ? _T_143 : 55'h0; // @[DivSqrtRecFN_small.scala 191:12]
  assign _T_145 = inReady & oddSqrt_S; // @[DivSqrtRecFN_small.scala 192:21]
  assign _T_149 = rawA_S_sig[52:51] - 2'h1; // @[DivSqrtRecFN_small.scala 193:56]
  assign _T_151 = {rawA_S_sig[50:0], 3'h0}; // @[DivSqrtRecFN_small.scala 194:44]
  assign _T_152 = {_T_149,_T_151}; // @[Cat.scala 30:58]
  assign _T_153 = _T_145 ? _T_152 : 56'h0; // @[DivSqrtRecFN_small.scala 192:12]
  assign _GEN_16 = {{1'd0}, _T_144}; // @[DivSqrtRecFN_small.scala 191:61]
  assign _T_154 = _GEN_16 | _T_153; // @[DivSqrtRecFN_small.scala 191:61]
  assign _T_156 = {rem_Z, 1'h0}; // @[DivSqrtRecFN_small.scala 198:29]
  assign _T_157 = inReady ? 56'h0 : _T_156; // @[DivSqrtRecFN_small.scala 198:12]
  assign rem = _T_154 | _T_157; // @[DivSqrtRecFN_small.scala 197:11]
  assign _T_158 = 64'h1 << cycleNum; // @[DivSqrtRecFN_small.scala 199:27]
  assign bitMask = _T_158[63:2]; // @[DivSqrtRecFN_small.scala 199:38]
  assign _T_160 = inReady & ~io_sqrtOp; // @[DivSqrtRecFN_small.scala 201:21]
  assign _T_161 = {rawB_S_sig, 1'h0}; // @[DivSqrtRecFN_small.scala 201:47]
  assign _T_162 = _T_160 ? _T_161 : 55'h0; // @[DivSqrtRecFN_small.scala 201:12]
  assign _T_163 = inReady & evenSqrt_S; // @[DivSqrtRecFN_small.scala 202:21]
  assign _T_164 = _T_163 ? 54'h20000000000000 : 54'h0; // @[DivSqrtRecFN_small.scala 202:12]
  assign _GEN_17 = {{1'd0}, _T_164}; // @[DivSqrtRecFN_small.scala 201:79]
  assign _T_165 = _T_162 | _GEN_17; // @[DivSqrtRecFN_small.scala 201:79]
  assign _T_167 = _T_145 ? 55'h50000000000000 : 55'h0; // @[DivSqrtRecFN_small.scala 203:12]
  assign _T_168 = _T_165 | _T_167; // @[DivSqrtRecFN_small.scala 202:79]
  assign _T_171 = ~inReady & ~sqrtOp_Z; // @[DivSqrtRecFN_small.scala 204:23]
  assign _T_172 = {1'h1,fractB_Z}; // @[Cat.scala 30:58]
  assign _T_173 = {_T_172, 1'h0}; // @[DivSqrtRecFN_small.scala 204:63]
  assign _T_174 = _T_171 ? _T_173 : 54'h0; // @[DivSqrtRecFN_small.scala 204:12]
  assign _GEN_18 = {{1'd0}, _T_174}; // @[DivSqrtRecFN_small.scala 203:79]
  assign _T_175 = _T_168 | _GEN_18; // @[DivSqrtRecFN_small.scala 203:79]
  assign _T_177 = ~inReady & sqrtOp_Z; // @[DivSqrtRecFN_small.scala 205:23]
  assign _T_178 = {sigX_Z, 1'h0}; // @[DivSqrtRecFN_small.scala 205:44]
  assign _GEN_19 = {{6'd0}, _T_178}; // @[DivSqrtRecFN_small.scala 205:48]
  assign _T_179 = _GEN_19 | bitMask; // @[DivSqrtRecFN_small.scala 205:48]
  assign _T_180 = _T_177 ? _T_179 : 62'h0; // @[DivSqrtRecFN_small.scala 205:12]
  assign _GEN_20 = {{7'd0}, _T_175}; // @[DivSqrtRecFN_small.scala 204:79]
  assign trialTerm = _GEN_20 | _T_180; // @[DivSqrtRecFN_small.scala 204:79]
  assign _T_181 = {1'b0,$signed(rem)}; // @[DivSqrtRecFN_small.scala 206:24]
  assign _T_182 = {1'b0,$signed(trialTerm)}; // @[DivSqrtRecFN_small.scala 206:41]
  assign _GEN_21 = {{6{_T_181[56]}},_T_181}; // @[DivSqrtRecFN_small.scala 206:29]
  assign trialRem = $signed(_GEN_21) - $signed(_T_182); // @[DivSqrtRecFN_small.scala 206:29]
  assign newBit = 63'sh0 <= $signed(trialRem); // @[DivSqrtRecFN_small.scala 207:27]
  assign _T_185 = cycleNum > 6'h2; // @[DivSqrtRecFN_small.scala 209:44]
  assign _T_186 = entering_normalCase | _T_185; // @[DivSqrtRecFN_small.scala 209:31]
  assign _T_187 = $signed(_GEN_21) - $signed(_T_182); // @[DivSqrtRecFN_small.scala 210:39]
  assign _T_188 = newBit ? _T_187 : {{7'd0}, rem}; // @[DivSqrtRecFN_small.scala 210:21]
  assign _GEN_10 = _T_186 ? _T_188 : {{8'd0}, rem_Z}; // @[DivSqrtRecFN_small.scala 209:56]
  assign _T_190 = ~inReady & newBit; // @[DivSqrtRecFN_small.scala 212:45]
  assign _T_191 = entering_normalCase | _T_190; // @[DivSqrtRecFN_small.scala 212:31]
  assign _T_192 = $signed(trialRem) != 63'sh0; // @[DivSqrtRecFN_small.scala 213:35]
  assign _T_195 = {newBit, 54'h0}; // @[DivSqrtRecFN_small.scala 215:47]
  assign _T_196 = _T_160 ? _T_195 : 55'h0; // @[DivSqrtRecFN_small.scala 215:16]
  assign _T_197 = inReady & io_sqrtOp; // @[DivSqrtRecFN_small.scala 216:25]
  assign _T_198 = _T_197 ? 54'h20000000000000 : 54'h0; // @[DivSqrtRecFN_small.scala 216:16]
  assign _GEN_22 = {{1'd0}, _T_198}; // @[DivSqrtRecFN_small.scala 215:77]
  assign _T_199 = _T_196 | _GEN_22; // @[DivSqrtRecFN_small.scala 215:77]
  assign _T_201 = {newBit, 52'h0}; // @[DivSqrtRecFN_small.scala 217:47]
  assign _T_202 = _T_145 ? _T_201 : 53'h0; // @[DivSqrtRecFN_small.scala 217:16]
  assign _GEN_23 = {{2'd0}, _T_202}; // @[DivSqrtRecFN_small.scala 216:77]
  assign _T_203 = _T_199 | _GEN_23; // @[DivSqrtRecFN_small.scala 216:77]
  assign _GEN_24 = {{7'd0}, sigX_Z}; // @[DivSqrtRecFN_small.scala 218:48]
  assign _T_205 = _GEN_24 | bitMask; // @[DivSqrtRecFN_small.scala 218:48]
  assign _T_206 = inReady ? 62'h0 : _T_205; // @[DivSqrtRecFN_small.scala 218:16]
  assign _GEN_25 = {{7'd0}, _T_203}; // @[DivSqrtRecFN_small.scala 217:77]
  assign _T_207 = _GEN_25 | _T_206; // @[DivSqrtRecFN_small.scala 217:77]
  assign _GEN_12 = _T_191 ? _T_207 : {{7'd0}, sigX_Z}; // @[DivSqrtRecFN_small.scala 212:57]
  assign rawOutValid = cycleNum == 6'h1; // @[DivSqrtRecFN_small.scala 223:33]
  assign _GEN_26 = {{55'd0}, notZeroRem_Z}; // @[DivSqrtRecFN_small.scala 235:35]
  assign io_inReady = cycleNum <= 6'h1; // @[DivSqrtRecFN_small.scala 164:16]
  assign io_rawOutValid_div = rawOutValid & ~sqrtOp_Z; // @[DivSqrtRecFN_small.scala 225:25]
  assign io_rawOutValid_sqrt = rawOutValid & sqrtOp_Z; // @[DivSqrtRecFN_small.scala 226:25]
  assign io_roundingModeOut = roundingMode_Z; // @[DivSqrtRecFN_small.scala 227:25]
  assign io_invalidExc = majorExc_Z & isNaN_Z; // @[DivSqrtRecFN_small.scala 228:22]
  assign io_infiniteExc = majorExc_Z & ~isNaN_Z; // @[DivSqrtRecFN_small.scala 229:22]
  assign io_rawOut_isNaN = isNaN_Z; // @[DivSqrtRecFN_small.scala 230:22]
  assign io_rawOut_isInf = isInf_Z; // @[DivSqrtRecFN_small.scala 231:22]
  assign io_rawOut_isZero = isZero_Z; // @[DivSqrtRecFN_small.scala 232:22]
  assign io_rawOut_sign = sign_Z; // @[DivSqrtRecFN_small.scala 233:22]
  assign io_rawOut_sExp = sExp_Z; // @[DivSqrtRecFN_small.scala 234:22]
  assign io_rawOut_sig = _T_178 | _GEN_26; // @[DivSqrtRecFN_small.scala 235:22]
  assign DivSqrtRecFNToRaw_small_1_cov_read_addr = DivSqrtRecFNToRaw_small_1_state;
  assign DivSqrtRecFNToRaw_small_1_cov_read_data = DivSqrtRecFNToRaw_small_1_cov[DivSqrtRecFNToRaw_small_1_cov_read_addr]; // @[Coverage map for DivSqrtRecFNToRaw_small_1]
  assign DivSqrtRecFNToRaw_small_1_cov_write_data = 1'h1;
  assign DivSqrtRecFNToRaw_small_1_cov_write_addr = DivSqrtRecFNToRaw_small_1_state;
  assign DivSqrtRecFNToRaw_small_1_cov_write_mask = 1'h1;
  assign DivSqrtRecFNToRaw_small_1_cov_write_en = 1'h1;
  assign sqrtOp_Z_shl = sqrtOp_Z;
  assign sqrtOp_Z_pad = {6'h0,sqrtOp_Z_shl};
  assign cycleNum_shl = {cycleNum, 1'h0};
  assign cycleNum_pad = cycleNum_shl;
  assign DivSqrtRecFNToRaw_small_1_xor0 = sqrtOp_Z_pad ^ cycleNum_pad;
  assign io_covSum = DivSqrtRecFNToRaw_small_1_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleNum = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sqrtOp_Z = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  majorExc_Z = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  isNaN_Z = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  isInf_Z = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  isZero_Z = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sign_Z = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  sExp_Z = _RAND_7[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {2{`RANDOM}};
  fractB_Z = _RAND_8[51:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  roundingMode_Z = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {2{`RANDOM}};
  rem_Z = _RAND_10[54:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  notZeroRem_Z = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {2{`RANDOM}};
  sigX_Z = _RAND_12[54:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  DivSqrtRecFNToRaw_small_1_state = _RAND_13[6:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    DivSqrtRecFNToRaw_small_1_cov[initvar] = _RAND_14[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  DivSqrtRecFNToRaw_small_1_covSum = _RAND_15[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      cycleNum <= 6'h0;
    end else if (reset) begin
      cycleNum <= 6'h0;
    end else if (_T_114) begin
      cycleNum <= _T_134;
    end
    if (metaReset) begin
      sqrtOp_Z <= 1'h0;
    end else if (entering) begin
      sqrtOp_Z <= io_sqrtOp;
    end
    if (metaReset) begin
      majorExc_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        majorExc_Z <= _T_71;
      end else begin
        majorExc_Z <= _T_84;
      end
    end
    if (metaReset) begin
      isNaN_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        isNaN_Z <= _T_85;
      end else begin
        isNaN_Z <= _T_87;
      end
    end
    if (metaReset) begin
      isInf_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        isInf_Z <= rawA_S_isInf;
      end else begin
        isInf_Z <= _T_88;
      end
    end
    if (metaReset) begin
      isZero_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        isZero_Z <= rawA_S_isZero;
      end else begin
        isZero_Z <= _T_89;
      end
    end
    if (metaReset) begin
      sign_Z <= 1'h0;
    end else if (entering) begin
      sign_Z <= sign_S;
    end
    if (metaReset) begin
      sExp_Z <= 13'h0;
    end else if (entering_normalCase) begin
      if (io_sqrtOp) begin
        sExp_Z <= _T_136;
      end else begin
        sExp_Z <= sSatExpQuot_S_div;
      end
    end
    if (metaReset) begin
      fractB_Z <= 52'h0;
    end else if (_T_139) begin
      fractB_Z <= rawB_S_sig[51:0];
    end
    if (metaReset) begin
      roundingMode_Z <= 3'h0;
    end else if (entering_normalCase) begin
      roundingMode_Z <= io_roundingMode;
    end
    if (metaReset) begin
      rem_Z <= 55'h0;
    end else begin
      rem_Z <= _GEN_10[54:0];
    end
    if (metaReset) begin
      notZeroRem_Z <= 1'h0;
    end else if (_T_191) begin
      notZeroRem_Z <= _T_192;
    end
    if (metaReset) begin
      sigX_Z <= 55'h0;
    end else begin
      sigX_Z <= _GEN_12[54:0];
    end
    DivSqrtRecFNToRaw_small_1_state <= DivSqrtRecFNToRaw_small_1_xor0;
    if (!(DivSqrtRecFNToRaw_small_1_cov_read_data)) begin
      DivSqrtRecFNToRaw_small_1_covSum <= DivSqrtRecFNToRaw_small_1_covSum + 1'h1;
    end
  end
  always @(posedge clock) begin
    if(DivSqrtRecFNToRaw_small_1_cov_write_en & DivSqrtRecFNToRaw_small_1_cov_write_mask) begin
      DivSqrtRecFNToRaw_small_1_cov[DivSqrtRecFNToRaw_small_1_cov_write_addr] <= DivSqrtRecFNToRaw_small_1_cov_write_data; // @[Coverage map for DivSqrtRecFNToRaw_small_1]
    end
  end
endmodule
module RoundRawFNToRecFN_3(
  input         io_invalidExc,
  input         io_infiniteExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [12:0] io_in_sExp,
  input  [55:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundAnyRawFNToRecFN_io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_infiniteExc; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [12:0] roundAnyRawFNToRecFN_io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [55:0] roundAnyRawFNToRecFN_io_in_sig; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [2:0] roundAnyRawFNToRecFN_io_roundingMode; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_detectTininess; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [64:0] roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [29:0] roundAnyRawFNToRecFN_io_covSum; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_metaAssert; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [29:0] RoundRawFNToRecFN_3_covSum;
  wire [29:0] roundAnyRawFNToRecFN_sum;
  wire  roundAnyRawFNToRecFN_metaAssert_wire;
  RoundAnyRawFNToRecFN_6 roundAnyRawFNToRecFN ( // @[RoundAnyRawFNToRecFN.scala 307:15]
    .io_invalidExc(roundAnyRawFNToRecFN_io_invalidExc),
    .io_infiniteExc(roundAnyRawFNToRecFN_io_infiniteExc),
    .io_in_isNaN(roundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundAnyRawFNToRecFN_io_detectTininess),
    .io_out(roundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundAnyRawFNToRecFN_io_covSum),
    .metaAssert(roundAnyRawFNToRecFN_metaAssert)
  );
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 315:23]
  assign io_exceptionFlags = roundAnyRawFNToRecFN_io_exceptionFlags; // @[RoundAnyRawFNToRecFN.scala 316:23]
  assign roundAnyRawFNToRecFN_io_invalidExc = io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 310:44]
  assign roundAnyRawFNToRecFN_io_infiniteExc = io_infiniteExc; // @[RoundAnyRawFNToRecFN.scala 311:44]
  assign roundAnyRawFNToRecFN_io_in_isNaN = io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isInf = io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isZero = io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_in_sign; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sig = io_in_sig; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[RoundAnyRawFNToRecFN.scala 313:44]
  assign roundAnyRawFNToRecFN_io_detectTininess = io_detectTininess; // @[RoundAnyRawFNToRecFN.scala 314:44]
  assign RoundRawFNToRecFN_3_covSum = 30'h0;
  assign roundAnyRawFNToRecFN_sum = RoundRawFNToRecFN_3_covSum + roundAnyRawFNToRecFN_io_covSum;
  assign io_covSum = roundAnyRawFNToRecFN_sum;
  assign roundAnyRawFNToRecFN_metaAssert_wire = roundAnyRawFNToRecFN_metaAssert;
  assign metaAssert = roundAnyRawFNToRecFN_metaAssert_wire;
endmodule
module RVCExpander(
  input  [31:0] io_in,
  output [31:0] io_out_bits,
  output [4:0]  io_out_rd,
  output [4:0]  io_out_rs1,
  output [4:0]  io_out_rs2,
  output [4:0]  io_out_rs3,
  output        io_rvc,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  _T_9; // @[RVC.scala 53:29]
  wire [6:0] _T_10; // @[RVC.scala 53:20]
  wire [4:0] _T_20; // @[Cat.scala 30:58]
  wire [29:0] _T_24; // @[Cat.scala 30:58]
  wire [7:0] _T_35; // @[Cat.scala 30:58]
  wire [4:0] _T_37; // @[Cat.scala 30:58]
  wire [27:0] _T_43; // @[Cat.scala 30:58]
  wire [6:0] _T_58; // @[Cat.scala 30:58]
  wire [26:0] _T_66; // @[Cat.scala 30:58]
  wire [27:0] _T_87; // @[Cat.scala 30:58]
  wire [26:0] _T_119; // @[Cat.scala 30:58]
  wire [27:0] _T_147; // @[Cat.scala 30:58]
  wire [26:0] _T_179; // @[Cat.scala 30:58]
  wire [27:0] _T_207; // @[Cat.scala 30:58]
  wire [6:0] _T_219; // @[Bitwise.scala 72:12]
  wire [11:0] _T_221; // @[Cat.scala 30:58]
  wire [31:0] _T_227; // @[Cat.scala 30:58]
  wire  _T_236; // @[RVC.scala 77:24]
  wire [6:0] _T_237; // @[RVC.scala 77:20]
  wire [31:0] _T_248; // @[Cat.scala 30:58]
  wire [31:0] _T_265; // @[Cat.scala 30:58]
  wire  _T_277; // @[RVC.scala 90:29]
  wire [6:0] _T_278; // @[RVC.scala 90:20]
  wire [14:0] _T_281; // @[Bitwise.scala 72:12]
  wire [31:0] _T_284; // @[Cat.scala 30:58]
  wire [31:0] _T_288; // @[Cat.scala 30:58]
  wire  _T_297; // @[RVC.scala 92:14]
  wire  _T_299; // @[RVC.scala 92:27]
  wire  _T_300; // @[RVC.scala 92:21]
  wire [6:0] _T_307; // @[RVC.scala 86:20]
  wire [2:0] _T_310; // @[Bitwise.scala 72:12]
  wire [31:0] _T_325; // @[Cat.scala 30:58]
  wire [31:0] _T_333_bits; // @[RVC.scala 92:10]
  wire [4:0] _T_333_rd; // @[RVC.scala 92:10]
  wire [4:0] _T_333_rs2; // @[RVC.scala 92:10]
  wire [4:0] _T_333_rs3; // @[RVC.scala 92:10]
  wire [25:0] _T_344; // @[Cat.scala 30:58]
  wire [30:0] _GEN_0; // @[RVC.scala 99:23]
  wire [30:0] _T_356; // @[RVC.scala 99:23]
  wire [31:0] _T_369; // @[Cat.scala 30:58]
  wire [2:0] _T_372; // @[Cat.scala 30:58]
  wire  _T_373; // @[package.scala 31:81]
  wire [2:0] _T_374; // @[package.scala 31:71]
  wire  _T_375; // @[package.scala 31:81]
  wire [2:0] _T_376; // @[package.scala 31:71]
  wire  _T_377; // @[package.scala 31:81]
  wire [2:0] _T_378; // @[package.scala 31:71]
  wire  _T_379; // @[package.scala 31:81]
  wire [2:0] _T_380; // @[package.scala 31:71]
  wire  _T_381; // @[package.scala 31:81]
  wire [2:0] _T_382; // @[package.scala 31:71]
  wire  _T_383; // @[package.scala 31:81]
  wire [2:0] _T_384; // @[package.scala 31:71]
  wire  _T_385; // @[package.scala 31:81]
  wire [2:0] _T_386; // @[package.scala 31:71]
  wire  _T_388; // @[RVC.scala 103:30]
  wire [30:0] _T_389; // @[RVC.scala 103:22]
  wire [6:0] _T_391; // @[RVC.scala 104:22]
  wire [24:0] _T_401; // @[Cat.scala 30:58]
  wire [30:0] _GEN_1; // @[RVC.scala 105:43]
  wire [30:0] _T_402; // @[RVC.scala 105:43]
  wire  _T_404; // @[package.scala 31:81]
  wire [30:0] _T_405; // @[package.scala 31:71]
  wire  _T_406; // @[package.scala 31:81]
  wire [31:0] _T_407; // @[package.scala 31:71]
  wire  _T_408; // @[package.scala 31:81]
  wire [31:0] _T_409; // @[package.scala 31:71]
  wire [9:0] _T_421; // @[Bitwise.scala 72:12]
  wire [20:0] _T_436; // @[Cat.scala 30:58]
  wire [31:0] _T_499; // @[Cat.scala 30:58]
  wire [4:0] _T_509; // @[Bitwise.scala 72:12]
  wire [12:0] _T_518; // @[Cat.scala 30:58]
  wire [31:0] _T_567; // @[Cat.scala 30:58]
  wire [31:0] _T_635; // @[Cat.scala 30:58]
  wire [6:0] _T_643; // @[RVC.scala 113:23]
  wire [25:0] _T_652; // @[Cat.scala 30:58]
  wire [28:0] _T_669; // @[Cat.scala 30:58]
  wire [27:0] _T_685; // @[Cat.scala 30:58]
  wire [28:0] _T_701; // @[Cat.scala 30:58]
  wire [24:0] _T_712; // @[Cat.scala 30:58]
  wire [24:0] _T_724; // @[Cat.scala 30:58]
  wire [24:0] _T_736; // @[Cat.scala 30:58]
  wire [24:0] _T_738; // @[Cat.scala 30:58]
  wire [24:0] _T_741; // @[RVC.scala 134:33]
  wire  _T_748; // @[RVC.scala 135:27]
  wire [31:0] _T_717_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _T_746_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _T_749_bits; // @[RVC.scala 135:22]
  wire [4:0] _T_749_rd; // @[RVC.scala 135:22]
  wire [4:0] _T_749_rs1; // @[RVC.scala 135:22]
  wire [4:0] _T_749_rs2; // @[RVC.scala 135:22]
  wire [4:0] _T_749_rs3; // @[RVC.scala 135:22]
  wire [24:0] _T_755; // @[Cat.scala 30:58]
  wire [24:0] _T_757; // @[Cat.scala 30:58]
  wire [24:0] _T_758; // @[RVC.scala 137:47]
  wire [24:0] _T_761; // @[RVC.scala 138:33]
  wire [31:0] _T_730_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _T_766_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _T_769_bits; // @[RVC.scala 139:25]
  wire [4:0] _T_769_rd; // @[RVC.scala 139:25]
  wire [4:0] _T_769_rs1; // @[RVC.scala 139:25]
  wire [31:0] _T_771_bits; // @[RVC.scala 140:10]
  wire [4:0] _T_771_rd; // @[RVC.scala 140:10]
  wire [4:0] _T_771_rs1; // @[RVC.scala 140:10]
  wire [4:0] _T_771_rs2; // @[RVC.scala 140:10]
  wire [4:0] _T_771_rs3; // @[RVC.scala 140:10]
  wire [8:0] _T_775; // @[Cat.scala 30:58]
  wire [28:0] _T_787; // @[Cat.scala 30:58]
  wire [7:0] _T_796; // @[Cat.scala 30:58]
  wire [27:0] _T_808; // @[Cat.scala 30:58]
  wire [28:0] _T_829; // @[Cat.scala 30:58]
  wire [4:0] _T_885; // @[Cat.scala 30:58]
  wire  _T_886; // @[package.scala 31:81]
  wire [31:0] _T_52_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _T_31_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _T_887_bits; // @[package.scala 31:71]
  wire [4:0] _T_887_rd; // @[package.scala 31:71]
  wire [4:0] _T_887_rs1; // @[package.scala 31:71]
  wire [4:0] _T_887_rs3; // @[package.scala 31:71]
  wire  _T_888; // @[package.scala 31:81]
  wire [31:0] _T_75_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _T_889_bits; // @[package.scala 31:71]
  wire [4:0] _T_889_rd; // @[package.scala 31:71]
  wire [4:0] _T_889_rs1; // @[package.scala 31:71]
  wire [4:0] _T_889_rs3; // @[package.scala 31:71]
  wire  _T_890; // @[package.scala 31:81]
  wire [31:0] _T_96_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _T_891_bits; // @[package.scala 31:71]
  wire [4:0] _T_891_rd; // @[package.scala 31:71]
  wire [4:0] _T_891_rs1; // @[package.scala 31:71]
  wire [4:0] _T_891_rs3; // @[package.scala 31:71]
  wire  _T_892; // @[package.scala 31:81]
  wire [31:0] _T_128_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _T_893_bits; // @[package.scala 31:71]
  wire [4:0] _T_893_rd; // @[package.scala 31:71]
  wire [4:0] _T_893_rs1; // @[package.scala 31:71]
  wire [4:0] _T_893_rs3; // @[package.scala 31:71]
  wire  _T_894; // @[package.scala 31:81]
  wire [31:0] _T_156_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _T_895_bits; // @[package.scala 31:71]
  wire [4:0] _T_895_rd; // @[package.scala 31:71]
  wire [4:0] _T_895_rs1; // @[package.scala 31:71]
  wire [4:0] _T_895_rs3; // @[package.scala 31:71]
  wire  _T_896; // @[package.scala 31:81]
  wire [31:0] _T_188_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _T_897_bits; // @[package.scala 31:71]
  wire [4:0] _T_897_rd; // @[package.scala 31:71]
  wire [4:0] _T_897_rs1; // @[package.scala 31:71]
  wire [4:0] _T_897_rs3; // @[package.scala 31:71]
  wire  _T_898; // @[package.scala 31:81]
  wire [31:0] _T_216_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _T_899_bits; // @[package.scala 31:71]
  wire [4:0] _T_899_rd; // @[package.scala 31:71]
  wire [4:0] _T_899_rs1; // @[package.scala 31:71]
  wire [4:0] _T_899_rs3; // @[package.scala 31:71]
  wire  _T_900; // @[package.scala 31:81]
  wire [31:0] _T_901_bits; // @[package.scala 31:71]
  wire [4:0] _T_901_rd; // @[package.scala 31:71]
  wire [4:0] _T_901_rs1; // @[package.scala 31:71]
  wire [4:0] _T_901_rs2; // @[package.scala 31:71]
  wire [4:0] _T_901_rs3; // @[package.scala 31:71]
  wire  _T_902; // @[package.scala 31:81]
  wire [31:0] _T_903_bits; // @[package.scala 31:71]
  wire [4:0] _T_903_rd; // @[package.scala 31:71]
  wire [4:0] _T_903_rs1; // @[package.scala 31:71]
  wire [4:0] _T_903_rs2; // @[package.scala 31:71]
  wire [4:0] _T_903_rs3; // @[package.scala 31:71]
  wire  _T_904; // @[package.scala 31:81]
  wire [31:0] _T_905_bits; // @[package.scala 31:71]
  wire [4:0] _T_905_rd; // @[package.scala 31:71]
  wire [4:0] _T_905_rs1; // @[package.scala 31:71]
  wire [4:0] _T_905_rs2; // @[package.scala 31:71]
  wire [4:0] _T_905_rs3; // @[package.scala 31:71]
  wire  _T_906; // @[package.scala 31:81]
  wire [31:0] _T_907_bits; // @[package.scala 31:71]
  wire [4:0] _T_907_rd; // @[package.scala 31:71]
  wire [4:0] _T_907_rs1; // @[package.scala 31:71]
  wire [4:0] _T_907_rs2; // @[package.scala 31:71]
  wire [4:0] _T_907_rs3; // @[package.scala 31:71]
  wire  _T_908; // @[package.scala 31:81]
  wire [31:0] _T_909_bits; // @[package.scala 31:71]
  wire [4:0] _T_909_rd; // @[package.scala 31:71]
  wire [4:0] _T_909_rs1; // @[package.scala 31:71]
  wire [4:0] _T_909_rs2; // @[package.scala 31:71]
  wire [4:0] _T_909_rs3; // @[package.scala 31:71]
  wire  _T_910; // @[package.scala 31:81]
  wire [31:0] _T_911_bits; // @[package.scala 31:71]
  wire [4:0] _T_911_rd; // @[package.scala 31:71]
  wire [4:0] _T_911_rs1; // @[package.scala 31:71]
  wire [4:0] _T_911_rs2; // @[package.scala 31:71]
  wire [4:0] _T_911_rs3; // @[package.scala 31:71]
  wire  _T_912; // @[package.scala 31:81]
  wire [31:0] _T_913_bits; // @[package.scala 31:71]
  wire [4:0] _T_913_rd; // @[package.scala 31:71]
  wire [4:0] _T_913_rs1; // @[package.scala 31:71]
  wire [4:0] _T_913_rs2; // @[package.scala 31:71]
  wire [4:0] _T_913_rs3; // @[package.scala 31:71]
  wire  _T_914; // @[package.scala 31:81]
  wire [31:0] _T_915_bits; // @[package.scala 31:71]
  wire [4:0] _T_915_rd; // @[package.scala 31:71]
  wire [4:0] _T_915_rs1; // @[package.scala 31:71]
  wire [4:0] _T_915_rs2; // @[package.scala 31:71]
  wire [4:0] _T_915_rs3; // @[package.scala 31:71]
  wire  _T_916; // @[package.scala 31:81]
  wire [31:0] _T_658_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _T_917_bits; // @[package.scala 31:71]
  wire [4:0] _T_917_rd; // @[package.scala 31:71]
  wire [4:0] _T_917_rs1; // @[package.scala 31:71]
  wire [4:0] _T_917_rs2; // @[package.scala 31:71]
  wire [4:0] _T_917_rs3; // @[package.scala 31:71]
  wire  _T_918; // @[package.scala 31:81]
  wire [31:0] _T_674_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _T_919_bits; // @[package.scala 31:71]
  wire [4:0] _T_919_rd; // @[package.scala 31:71]
  wire [4:0] _T_919_rs1; // @[package.scala 31:71]
  wire [4:0] _T_919_rs2; // @[package.scala 31:71]
  wire [4:0] _T_919_rs3; // @[package.scala 31:71]
  wire  _T_920; // @[package.scala 31:81]
  wire [31:0] _T_690_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _T_921_bits; // @[package.scala 31:71]
  wire [4:0] _T_921_rd; // @[package.scala 31:71]
  wire [4:0] _T_921_rs1; // @[package.scala 31:71]
  wire [4:0] _T_921_rs2; // @[package.scala 31:71]
  wire [4:0] _T_921_rs3; // @[package.scala 31:71]
  wire  _T_922; // @[package.scala 31:81]
  wire [31:0] _T_706_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _T_923_bits; // @[package.scala 31:71]
  wire [4:0] _T_923_rd; // @[package.scala 31:71]
  wire [4:0] _T_923_rs1; // @[package.scala 31:71]
  wire [4:0] _T_923_rs2; // @[package.scala 31:71]
  wire [4:0] _T_923_rs3; // @[package.scala 31:71]
  wire  _T_924; // @[package.scala 31:81]
  wire [31:0] _T_925_bits; // @[package.scala 31:71]
  wire [4:0] _T_925_rd; // @[package.scala 31:71]
  wire [4:0] _T_925_rs1; // @[package.scala 31:71]
  wire [4:0] _T_925_rs2; // @[package.scala 31:71]
  wire [4:0] _T_925_rs3; // @[package.scala 31:71]
  wire  _T_926; // @[package.scala 31:81]
  wire [31:0] _T_792_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _T_927_bits; // @[package.scala 31:71]
  wire [4:0] _T_927_rd; // @[package.scala 31:71]
  wire [4:0] _T_927_rs1; // @[package.scala 31:71]
  wire [4:0] _T_927_rs2; // @[package.scala 31:71]
  wire [4:0] _T_927_rs3; // @[package.scala 31:71]
  wire  _T_928; // @[package.scala 31:81]
  wire [31:0] _T_813_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _T_929_bits; // @[package.scala 31:71]
  wire [4:0] _T_929_rd; // @[package.scala 31:71]
  wire [4:0] _T_929_rs1; // @[package.scala 31:71]
  wire [4:0] _T_929_rs2; // @[package.scala 31:71]
  wire [4:0] _T_929_rs3; // @[package.scala 31:71]
  wire  _T_930; // @[package.scala 31:81]
  wire [31:0] _T_834_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _T_931_bits; // @[package.scala 31:71]
  wire [4:0] _T_931_rd; // @[package.scala 31:71]
  wire [4:0] _T_931_rs1; // @[package.scala 31:71]
  wire [4:0] _T_931_rs2; // @[package.scala 31:71]
  wire [4:0] _T_931_rs3; // @[package.scala 31:71]
  wire  _T_932; // @[package.scala 31:81]
  wire [31:0] _T_933_bits; // @[package.scala 31:71]
  wire [4:0] _T_933_rd; // @[package.scala 31:71]
  wire [4:0] _T_933_rs1; // @[package.scala 31:71]
  wire [4:0] _T_933_rs2; // @[package.scala 31:71]
  wire [4:0] _T_933_rs3; // @[package.scala 31:71]
  wire  _T_934; // @[package.scala 31:81]
  wire [31:0] _T_935_bits; // @[package.scala 31:71]
  wire [4:0] _T_935_rd; // @[package.scala 31:71]
  wire [4:0] _T_935_rs1; // @[package.scala 31:71]
  wire [4:0] _T_935_rs2; // @[package.scala 31:71]
  wire [4:0] _T_935_rs3; // @[package.scala 31:71]
  wire  _T_936; // @[package.scala 31:81]
  wire [31:0] _T_937_bits; // @[package.scala 31:71]
  wire [4:0] _T_937_rd; // @[package.scala 31:71]
  wire [4:0] _T_937_rs1; // @[package.scala 31:71]
  wire [4:0] _T_937_rs2; // @[package.scala 31:71]
  wire [4:0] _T_937_rs3; // @[package.scala 31:71]
  wire  _T_938; // @[package.scala 31:81]
  wire [31:0] _T_939_bits; // @[package.scala 31:71]
  wire [4:0] _T_939_rd; // @[package.scala 31:71]
  wire [4:0] _T_939_rs1; // @[package.scala 31:71]
  wire [4:0] _T_939_rs2; // @[package.scala 31:71]
  wire [4:0] _T_939_rs3; // @[package.scala 31:71]
  wire  _T_940; // @[package.scala 31:81]
  wire [31:0] _T_941_bits; // @[package.scala 31:71]
  wire [4:0] _T_941_rd; // @[package.scala 31:71]
  wire [4:0] _T_941_rs1; // @[package.scala 31:71]
  wire [4:0] _T_941_rs2; // @[package.scala 31:71]
  wire [4:0] _T_941_rs3; // @[package.scala 31:71]
  wire  _T_942; // @[package.scala 31:81]
  wire [31:0] _T_943_bits; // @[package.scala 31:71]
  wire [4:0] _T_943_rd; // @[package.scala 31:71]
  wire [4:0] _T_943_rs1; // @[package.scala 31:71]
  wire [4:0] _T_943_rs2; // @[package.scala 31:71]
  wire [4:0] _T_943_rs3; // @[package.scala 31:71]
  wire  _T_944; // @[package.scala 31:81]
  wire [31:0] _T_945_bits; // @[package.scala 31:71]
  wire [4:0] _T_945_rd; // @[package.scala 31:71]
  wire [4:0] _T_945_rs1; // @[package.scala 31:71]
  wire [4:0] _T_945_rs2; // @[package.scala 31:71]
  wire [4:0] _T_945_rs3; // @[package.scala 31:71]
  wire  _T_946; // @[package.scala 31:81]
  wire [29:0] RVCExpander_covSum;
  assign _T_9 = io_in[12:5] != 8'h0; // @[RVC.scala 53:29]
  assign _T_10 = _T_9 ? 7'h13 : 7'h1f; // @[RVC.scala 53:20]
  assign _T_20 = {2'h1,io_in[4:2]}; // @[Cat.scala 30:58]
  assign _T_24 = {io_in[10:7],io_in[12:11],io_in[5],io_in[6],2'h0,5'h2,3'h0,2'h1,io_in[4:2],_T_10}; // @[Cat.scala 30:58]
  assign _T_35 = {io_in[6:5],io_in[12:10],3'h0}; // @[Cat.scala 30:58]
  assign _T_37 = {2'h1,io_in[9:7]}; // @[Cat.scala 30:58]
  assign _T_43 = {io_in[6:5],io_in[12:10],3'h0,2'h1,io_in[9:7],3'h3,2'h1,io_in[4:2],7'h7}; // @[Cat.scala 30:58]
  assign _T_58 = {io_in[5],io_in[12:10],io_in[6],2'h0}; // @[Cat.scala 30:58]
  assign _T_66 = {io_in[5],io_in[12:10],io_in[6],2'h0,2'h1,io_in[9:7],3'h2,2'h1,io_in[4:2],7'h3}; // @[Cat.scala 30:58]
  assign _T_87 = {io_in[6:5],io_in[12:10],3'h0,2'h1,io_in[9:7],3'h3,2'h1,io_in[4:2],7'h3}; // @[Cat.scala 30:58]
  assign _T_119 = {_T_58[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_T_58[4:0],7'h3f}; // @[Cat.scala 30:58]
  assign _T_147 = {_T_35[7:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,_T_35[4:0],7'h27}; // @[Cat.scala 30:58]
  assign _T_179 = {_T_58[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_T_58[4:0],7'h23}; // @[Cat.scala 30:58]
  assign _T_207 = {_T_35[7:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,_T_35[4:0],7'h23}; // @[Cat.scala 30:58]
  assign _T_219 = io_in[12] ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12]
  assign _T_221 = {_T_219,io_in[6:2]}; // @[Cat.scala 30:58]
  assign _T_227 = {_T_219,io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h13}; // @[Cat.scala 30:58]
  assign _T_236 = io_in[11:7] != 5'h0; // @[RVC.scala 77:24]
  assign _T_237 = _T_236 ? 7'h1b : 7'h1f; // @[RVC.scala 77:20]
  assign _T_248 = {_T_219,io_in[6:2],io_in[11:7],3'h0,io_in[11:7],_T_237}; // @[Cat.scala 30:58]
  assign _T_265 = {_T_219,io_in[6:2],5'h0,3'h0,io_in[11:7],7'h13}; // @[Cat.scala 30:58]
  assign _T_277 = _T_221 != 12'h0; // @[RVC.scala 90:29]
  assign _T_278 = _T_277 ? 7'h37 : 7'h3f; // @[RVC.scala 90:20]
  assign _T_281 = io_in[12] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  assign _T_284 = {_T_281,io_in[6:2],12'h0}; // @[Cat.scala 30:58]
  assign _T_288 = {_T_284[31:12],io_in[11:7],_T_278}; // @[Cat.scala 30:58]
  assign _T_297 = io_in[11:7] == 5'h0; // @[RVC.scala 92:14]
  assign _T_299 = io_in[11:7] == 5'h2; // @[RVC.scala 92:27]
  assign _T_300 = _T_297 | _T_299; // @[RVC.scala 92:21]
  assign _T_307 = _T_277 ? 7'h13 : 7'h1f; // @[RVC.scala 86:20]
  assign _T_310 = io_in[12] ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  assign _T_325 = {_T_310,io_in[4:3],io_in[5],io_in[2],io_in[6],4'h0,io_in[11:7],3'h0,io_in[11:7],_T_307}; // @[Cat.scala 30:58]
  assign _T_333_bits = _T_300 ? _T_325 : _T_288; // @[RVC.scala 92:10]
  assign _T_333_rd = _T_300 ? io_in[11:7] : io_in[11:7]; // @[RVC.scala 92:10]
  assign _T_333_rs2 = _T_300 ? _T_20 : _T_20; // @[RVC.scala 92:10]
  assign _T_333_rs3 = _T_300 ? io_in[31:27] : io_in[31:27]; // @[RVC.scala 92:10]
  assign _T_344 = {io_in[12],io_in[6:2],2'h1,io_in[9:7],3'h5,2'h1,io_in[9:7],7'h13}; // @[Cat.scala 30:58]
  assign _GEN_0 = {{5'd0}, _T_344}; // @[RVC.scala 99:23]
  assign _T_356 = _GEN_0 | 31'h40000000; // @[RVC.scala 99:23]
  assign _T_369 = {_T_219,io_in[6:2],2'h1,io_in[9:7],3'h7,2'h1,io_in[9:7],7'h13}; // @[Cat.scala 30:58]
  assign _T_372 = {io_in[12],io_in[6:5]}; // @[Cat.scala 30:58]
  assign _T_373 = _T_372 == 3'h1; // @[package.scala 31:81]
  assign _T_374 = _T_373 ? 3'h4 : 3'h0; // @[package.scala 31:71]
  assign _T_375 = _T_372 == 3'h2; // @[package.scala 31:81]
  assign _T_376 = _T_375 ? 3'h6 : _T_374; // @[package.scala 31:71]
  assign _T_377 = _T_372 == 3'h3; // @[package.scala 31:81]
  assign _T_378 = _T_377 ? 3'h7 : _T_376; // @[package.scala 31:71]
  assign _T_379 = _T_372 == 3'h4; // @[package.scala 31:81]
  assign _T_380 = _T_379 ? 3'h0 : _T_378; // @[package.scala 31:71]
  assign _T_381 = _T_372 == 3'h5; // @[package.scala 31:81]
  assign _T_382 = _T_381 ? 3'h0 : _T_380; // @[package.scala 31:71]
  assign _T_383 = _T_372 == 3'h6; // @[package.scala 31:81]
  assign _T_384 = _T_383 ? 3'h2 : _T_382; // @[package.scala 31:71]
  assign _T_385 = _T_372 == 3'h7; // @[package.scala 31:81]
  assign _T_386 = _T_385 ? 3'h3 : _T_384; // @[package.scala 31:71]
  assign _T_388 = io_in[6:5] == 2'h0; // @[RVC.scala 103:30]
  assign _T_389 = _T_388 ? 31'h40000000 : 31'h0; // @[RVC.scala 103:22]
  assign _T_391 = io_in[12] ? 7'h3b : 7'h33; // @[RVC.scala 104:22]
  assign _T_401 = {2'h1,io_in[4:2],2'h1,io_in[9:7],_T_386,2'h1,io_in[9:7],_T_391}; // @[Cat.scala 30:58]
  assign _GEN_1 = {{6'd0}, _T_401}; // @[RVC.scala 105:43]
  assign _T_402 = _GEN_1 | _T_389; // @[RVC.scala 105:43]
  assign _T_404 = io_in[11:10] == 2'h1; // @[package.scala 31:81]
  assign _T_405 = _T_404 ? _T_356 : {{5'd0}, _T_344}; // @[package.scala 31:71]
  assign _T_406 = io_in[11:10] == 2'h2; // @[package.scala 31:81]
  assign _T_407 = _T_406 ? _T_369 : {{1'd0}, _T_405}; // @[package.scala 31:71]
  assign _T_408 = io_in[11:10] == 2'h3; // @[package.scala 31:81]
  assign _T_409 = _T_408 ? {{1'd0}, _T_402} : _T_407; // @[package.scala 31:71]
  assign _T_421 = io_in[12] ? 10'h3ff : 10'h0; // @[Bitwise.scala 72:12]
  assign _T_436 = {_T_421,io_in[8],io_in[10:9],io_in[6],io_in[7],io_in[2],io_in[11],io_in[5:3],1'h0}; // @[Cat.scala 30:58]
  assign _T_499 = {_T_436[20],_T_436[10:1],_T_436[11],_T_436[19:12],5'h0,7'h6f}; // @[Cat.scala 30:58]
  assign _T_509 = io_in[12] ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12]
  assign _T_518 = {_T_509,io_in[6:5],io_in[2],io_in[11:10],io_in[4:3],1'h0}; // @[Cat.scala 30:58]
  assign _T_567 = {_T_518[12],_T_518[10:5],5'h0,2'h1,io_in[9:7],3'h0,_T_518[4:1],_T_518[11],7'h63}; // @[Cat.scala 30:58]
  assign _T_635 = {_T_518[12],_T_518[10:5],5'h0,2'h1,io_in[9:7],3'h1,_T_518[4:1],_T_518[11],7'h63}; // @[Cat.scala 30:58]
  assign _T_643 = _T_236 ? 7'h3 : 7'h1f; // @[RVC.scala 113:23]
  assign _T_652 = {io_in[12],io_in[6:2],io_in[11:7],3'h1,io_in[11:7],7'h13}; // @[Cat.scala 30:58]
  assign _T_669 = {io_in[4:2],io_in[12],io_in[6:5],3'h0,5'h2,3'h3,io_in[11:7],7'h7}; // @[Cat.scala 30:58]
  assign _T_685 = {io_in[3:2],io_in[12],io_in[6:4],2'h0,5'h2,3'h2,io_in[11:7],_T_643}; // @[Cat.scala 30:58]
  assign _T_701 = {io_in[4:2],io_in[12],io_in[6:5],3'h0,5'h2,3'h3,io_in[11:7],_T_643}; // @[Cat.scala 30:58]
  assign _T_712 = {io_in[6:2],5'h0,3'h0,io_in[11:7],7'h33}; // @[Cat.scala 30:58]
  assign _T_724 = {io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h33}; // @[Cat.scala 30:58]
  assign _T_736 = {io_in[6:2],io_in[11:7],3'h0,12'h67}; // @[Cat.scala 30:58]
  assign _T_738 = {_T_736[24:7],7'h1f}; // @[Cat.scala 30:58]
  assign _T_741 = _T_236 ? _T_736 : _T_738; // @[RVC.scala 134:33]
  assign _T_748 = io_in[6:2] != 5'h0; // @[RVC.scala 135:27]
  assign _T_717_bits = {{7'd0}, _T_712}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _T_746_bits = {{7'd0}, _T_741}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _T_749_bits = _T_748 ? _T_717_bits : _T_746_bits; // @[RVC.scala 135:22]
  assign _T_749_rd = _T_748 ? io_in[11:7] : 5'h0; // @[RVC.scala 135:22]
  assign _T_749_rs1 = _T_748 ? 5'h0 : io_in[11:7]; // @[RVC.scala 135:22]
  assign _T_749_rs2 = _T_748 ? io_in[6:2] : io_in[6:2]; // @[RVC.scala 135:22]
  assign _T_749_rs3 = _T_748 ? io_in[31:27] : io_in[31:27]; // @[RVC.scala 135:22]
  assign _T_755 = {io_in[6:2],io_in[11:7],3'h0,12'he7}; // @[Cat.scala 30:58]
  assign _T_757 = {_T_736[24:7],7'h73}; // @[Cat.scala 30:58]
  assign _T_758 = _T_757 | 25'h100000; // @[RVC.scala 137:47]
  assign _T_761 = _T_236 ? _T_755 : _T_758; // @[RVC.scala 138:33]
  assign _T_730_bits = {{7'd0}, _T_724}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _T_766_bits = {{7'd0}, _T_761}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _T_769_bits = _T_748 ? _T_730_bits : _T_766_bits; // @[RVC.scala 139:25]
  assign _T_769_rd = _T_748 ? io_in[11:7] : 5'h1; // @[RVC.scala 139:25]
  assign _T_769_rs1 = _T_748 ? io_in[11:7] : io_in[11:7]; // @[RVC.scala 139:25]
  assign _T_771_bits = io_in[12] ? _T_769_bits : _T_749_bits; // @[RVC.scala 140:10]
  assign _T_771_rd = io_in[12] ? _T_769_rd : _T_749_rd; // @[RVC.scala 140:10]
  assign _T_771_rs1 = io_in[12] ? _T_769_rs1 : _T_749_rs1; // @[RVC.scala 140:10]
  assign _T_771_rs2 = io_in[12] ? _T_749_rs2 : _T_749_rs2; // @[RVC.scala 140:10]
  assign _T_771_rs3 = io_in[12] ? _T_749_rs3 : _T_749_rs3; // @[RVC.scala 140:10]
  assign _T_775 = {io_in[9:7],io_in[12:10],3'h0}; // @[Cat.scala 30:58]
  assign _T_787 = {_T_775[8:5],io_in[6:2],5'h2,3'h3,_T_775[4:0],7'h27}; // @[Cat.scala 30:58]
  assign _T_796 = {io_in[8:7],io_in[12:9],2'h0}; // @[Cat.scala 30:58]
  assign _T_808 = {_T_796[7:5],io_in[6:2],5'h2,3'h2,_T_796[4:0],7'h23}; // @[Cat.scala 30:58]
  assign _T_829 = {_T_775[8:5],io_in[6:2],5'h2,3'h3,_T_775[4:0],7'h23}; // @[Cat.scala 30:58]
  assign _T_885 = {io_in[1:0],io_in[15:13]}; // @[Cat.scala 30:58]
  assign _T_886 = _T_885 == 5'h1; // @[package.scala 31:81]
  assign _T_52_bits = {{4'd0}, _T_43}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _T_31_bits = {{2'd0}, _T_24}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _T_887_bits = _T_886 ? _T_52_bits : _T_31_bits; // @[package.scala 31:71]
  assign _T_887_rd = _T_886 ? _T_20 : _T_20; // @[package.scala 31:71]
  assign _T_887_rs1 = _T_886 ? _T_37 : 5'h2; // @[package.scala 31:71]
  assign _T_887_rs3 = _T_886 ? io_in[31:27] : io_in[31:27]; // @[package.scala 31:71]
  assign _T_888 = _T_885 == 5'h2; // @[package.scala 31:81]
  assign _T_75_bits = {{5'd0}, _T_66}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _T_889_bits = _T_888 ? _T_75_bits : _T_887_bits; // @[package.scala 31:71]
  assign _T_889_rd = _T_888 ? _T_20 : _T_887_rd; // @[package.scala 31:71]
  assign _T_889_rs1 = _T_888 ? _T_37 : _T_887_rs1; // @[package.scala 31:71]
  assign _T_889_rs3 = _T_888 ? io_in[31:27] : _T_887_rs3; // @[package.scala 31:71]
  assign _T_890 = _T_885 == 5'h3; // @[package.scala 31:81]
  assign _T_96_bits = {{4'd0}, _T_87}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _T_891_bits = _T_890 ? _T_96_bits : _T_889_bits; // @[package.scala 31:71]
  assign _T_891_rd = _T_890 ? _T_20 : _T_889_rd; // @[package.scala 31:71]
  assign _T_891_rs1 = _T_890 ? _T_37 : _T_889_rs1; // @[package.scala 31:71]
  assign _T_891_rs3 = _T_890 ? io_in[31:27] : _T_889_rs3; // @[package.scala 31:71]
  assign _T_892 = _T_885 == 5'h4; // @[package.scala 31:81]
  assign _T_128_bits = {{5'd0}, _T_119}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _T_893_bits = _T_892 ? _T_128_bits : _T_891_bits; // @[package.scala 31:71]
  assign _T_893_rd = _T_892 ? _T_20 : _T_891_rd; // @[package.scala 31:71]
  assign _T_893_rs1 = _T_892 ? _T_37 : _T_891_rs1; // @[package.scala 31:71]
  assign _T_893_rs3 = _T_892 ? io_in[31:27] : _T_891_rs3; // @[package.scala 31:71]
  assign _T_894 = _T_885 == 5'h5; // @[package.scala 31:81]
  assign _T_156_bits = {{4'd0}, _T_147}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _T_895_bits = _T_894 ? _T_156_bits : _T_893_bits; // @[package.scala 31:71]
  assign _T_895_rd = _T_894 ? _T_20 : _T_893_rd; // @[package.scala 31:71]
  assign _T_895_rs1 = _T_894 ? _T_37 : _T_893_rs1; // @[package.scala 31:71]
  assign _T_895_rs3 = _T_894 ? io_in[31:27] : _T_893_rs3; // @[package.scala 31:71]
  assign _T_896 = _T_885 == 5'h6; // @[package.scala 31:81]
  assign _T_188_bits = {{5'd0}, _T_179}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _T_897_bits = _T_896 ? _T_188_bits : _T_895_bits; // @[package.scala 31:71]
  assign _T_897_rd = _T_896 ? _T_20 : _T_895_rd; // @[package.scala 31:71]
  assign _T_897_rs1 = _T_896 ? _T_37 : _T_895_rs1; // @[package.scala 31:71]
  assign _T_897_rs3 = _T_896 ? io_in[31:27] : _T_895_rs3; // @[package.scala 31:71]
  assign _T_898 = _T_885 == 5'h7; // @[package.scala 31:81]
  assign _T_216_bits = {{4'd0}, _T_207}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _T_899_bits = _T_898 ? _T_216_bits : _T_897_bits; // @[package.scala 31:71]
  assign _T_899_rd = _T_898 ? _T_20 : _T_897_rd; // @[package.scala 31:71]
  assign _T_899_rs1 = _T_898 ? _T_37 : _T_897_rs1; // @[package.scala 31:71]
  assign _T_899_rs3 = _T_898 ? io_in[31:27] : _T_897_rs3; // @[package.scala 31:71]
  assign _T_900 = _T_885 == 5'h8; // @[package.scala 31:81]
  assign _T_901_bits = _T_900 ? _T_227 : _T_899_bits; // @[package.scala 31:71]
  assign _T_901_rd = _T_900 ? io_in[11:7] : _T_899_rd; // @[package.scala 31:71]
  assign _T_901_rs1 = _T_900 ? io_in[11:7] : _T_899_rs1; // @[package.scala 31:71]
  assign _T_901_rs2 = _T_900 ? _T_20 : _T_899_rd; // @[package.scala 31:71]
  assign _T_901_rs3 = _T_900 ? io_in[31:27] : _T_899_rs3; // @[package.scala 31:71]
  assign _T_902 = _T_885 == 5'h9; // @[package.scala 31:81]
  assign _T_903_bits = _T_902 ? _T_248 : _T_901_bits; // @[package.scala 31:71]
  assign _T_903_rd = _T_902 ? io_in[11:7] : _T_901_rd; // @[package.scala 31:71]
  assign _T_903_rs1 = _T_902 ? io_in[11:7] : _T_901_rs1; // @[package.scala 31:71]
  assign _T_903_rs2 = _T_902 ? _T_20 : _T_901_rs2; // @[package.scala 31:71]
  assign _T_903_rs3 = _T_902 ? io_in[31:27] : _T_901_rs3; // @[package.scala 31:71]
  assign _T_904 = _T_885 == 5'ha; // @[package.scala 31:81]
  assign _T_905_bits = _T_904 ? _T_265 : _T_903_bits; // @[package.scala 31:71]
  assign _T_905_rd = _T_904 ? io_in[11:7] : _T_903_rd; // @[package.scala 31:71]
  assign _T_905_rs1 = _T_904 ? 5'h0 : _T_903_rs1; // @[package.scala 31:71]
  assign _T_905_rs2 = _T_904 ? _T_20 : _T_903_rs2; // @[package.scala 31:71]
  assign _T_905_rs3 = _T_904 ? io_in[31:27] : _T_903_rs3; // @[package.scala 31:71]
  assign _T_906 = _T_885 == 5'hb; // @[package.scala 31:81]
  assign _T_907_bits = _T_906 ? _T_333_bits : _T_905_bits; // @[package.scala 31:71]
  assign _T_907_rd = _T_906 ? _T_333_rd : _T_905_rd; // @[package.scala 31:71]
  assign _T_907_rs1 = _T_906 ? _T_333_rd : _T_905_rs1; // @[package.scala 31:71]
  assign _T_907_rs2 = _T_906 ? _T_333_rs2 : _T_905_rs2; // @[package.scala 31:71]
  assign _T_907_rs3 = _T_906 ? _T_333_rs3 : _T_905_rs3; // @[package.scala 31:71]
  assign _T_908 = _T_885 == 5'hc; // @[package.scala 31:81]
  assign _T_909_bits = _T_908 ? _T_409 : _T_907_bits; // @[package.scala 31:71]
  assign _T_909_rd = _T_908 ? _T_37 : _T_907_rd; // @[package.scala 31:71]
  assign _T_909_rs1 = _T_908 ? _T_37 : _T_907_rs1; // @[package.scala 31:71]
  assign _T_909_rs2 = _T_908 ? _T_20 : _T_907_rs2; // @[package.scala 31:71]
  assign _T_909_rs3 = _T_908 ? io_in[31:27] : _T_907_rs3; // @[package.scala 31:71]
  assign _T_910 = _T_885 == 5'hd; // @[package.scala 31:81]
  assign _T_911_bits = _T_910 ? _T_499 : _T_909_bits; // @[package.scala 31:71]
  assign _T_911_rd = _T_910 ? 5'h0 : _T_909_rd; // @[package.scala 31:71]
  assign _T_911_rs1 = _T_910 ? _T_37 : _T_909_rs1; // @[package.scala 31:71]
  assign _T_911_rs2 = _T_910 ? _T_20 : _T_909_rs2; // @[package.scala 31:71]
  assign _T_911_rs3 = _T_910 ? io_in[31:27] : _T_909_rs3; // @[package.scala 31:71]
  assign _T_912 = _T_885 == 5'he; // @[package.scala 31:81]
  assign _T_913_bits = _T_912 ? _T_567 : _T_911_bits; // @[package.scala 31:71]
  assign _T_913_rd = _T_912 ? _T_37 : _T_911_rd; // @[package.scala 31:71]
  assign _T_913_rs1 = _T_912 ? _T_37 : _T_911_rs1; // @[package.scala 31:71]
  assign _T_913_rs2 = _T_912 ? 5'h0 : _T_911_rs2; // @[package.scala 31:71]
  assign _T_913_rs3 = _T_912 ? io_in[31:27] : _T_911_rs3; // @[package.scala 31:71]
  assign _T_914 = _T_885 == 5'hf; // @[package.scala 31:81]
  assign _T_915_bits = _T_914 ? _T_635 : _T_913_bits; // @[package.scala 31:71]
  assign _T_915_rd = _T_914 ? 5'h0 : _T_913_rd; // @[package.scala 31:71]
  assign _T_915_rs1 = _T_914 ? _T_37 : _T_913_rs1; // @[package.scala 31:71]
  assign _T_915_rs2 = _T_914 ? 5'h0 : _T_913_rs2; // @[package.scala 31:71]
  assign _T_915_rs3 = _T_914 ? io_in[31:27] : _T_913_rs3; // @[package.scala 31:71]
  assign _T_916 = _T_885 == 5'h10; // @[package.scala 31:81]
  assign _T_658_bits = {{6'd0}, _T_652}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _T_917_bits = _T_916 ? _T_658_bits : _T_915_bits; // @[package.scala 31:71]
  assign _T_917_rd = _T_916 ? io_in[11:7] : _T_915_rd; // @[package.scala 31:71]
  assign _T_917_rs1 = _T_916 ? io_in[11:7] : _T_915_rs1; // @[package.scala 31:71]
  assign _T_917_rs2 = _T_916 ? io_in[6:2] : _T_915_rs2; // @[package.scala 31:71]
  assign _T_917_rs3 = _T_916 ? io_in[31:27] : _T_915_rs3; // @[package.scala 31:71]
  assign _T_918 = _T_885 == 5'h11; // @[package.scala 31:81]
  assign _T_674_bits = {{3'd0}, _T_669}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _T_919_bits = _T_918 ? _T_674_bits : _T_917_bits; // @[package.scala 31:71]
  assign _T_919_rd = _T_918 ? io_in[11:7] : _T_917_rd; // @[package.scala 31:71]
  assign _T_919_rs1 = _T_918 ? 5'h2 : _T_917_rs1; // @[package.scala 31:71]
  assign _T_919_rs2 = _T_918 ? io_in[6:2] : _T_917_rs2; // @[package.scala 31:71]
  assign _T_919_rs3 = _T_918 ? io_in[31:27] : _T_917_rs3; // @[package.scala 31:71]
  assign _T_920 = _T_885 == 5'h12; // @[package.scala 31:81]
  assign _T_690_bits = {{4'd0}, _T_685}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _T_921_bits = _T_920 ? _T_690_bits : _T_919_bits; // @[package.scala 31:71]
  assign _T_921_rd = _T_920 ? io_in[11:7] : _T_919_rd; // @[package.scala 31:71]
  assign _T_921_rs1 = _T_920 ? 5'h2 : _T_919_rs1; // @[package.scala 31:71]
  assign _T_921_rs2 = _T_920 ? io_in[6:2] : _T_919_rs2; // @[package.scala 31:71]
  assign _T_921_rs3 = _T_920 ? io_in[31:27] : _T_919_rs3; // @[package.scala 31:71]
  assign _T_922 = _T_885 == 5'h13; // @[package.scala 31:81]
  assign _T_706_bits = {{3'd0}, _T_701}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _T_923_bits = _T_922 ? _T_706_bits : _T_921_bits; // @[package.scala 31:71]
  assign _T_923_rd = _T_922 ? io_in[11:7] : _T_921_rd; // @[package.scala 31:71]
  assign _T_923_rs1 = _T_922 ? 5'h2 : _T_921_rs1; // @[package.scala 31:71]
  assign _T_923_rs2 = _T_922 ? io_in[6:2] : _T_921_rs2; // @[package.scala 31:71]
  assign _T_923_rs3 = _T_922 ? io_in[31:27] : _T_921_rs3; // @[package.scala 31:71]
  assign _T_924 = _T_885 == 5'h14; // @[package.scala 31:81]
  assign _T_925_bits = _T_924 ? _T_771_bits : _T_923_bits; // @[package.scala 31:71]
  assign _T_925_rd = _T_924 ? _T_771_rd : _T_923_rd; // @[package.scala 31:71]
  assign _T_925_rs1 = _T_924 ? _T_771_rs1 : _T_923_rs1; // @[package.scala 31:71]
  assign _T_925_rs2 = _T_924 ? _T_771_rs2 : _T_923_rs2; // @[package.scala 31:71]
  assign _T_925_rs3 = _T_924 ? _T_771_rs3 : _T_923_rs3; // @[package.scala 31:71]
  assign _T_926 = _T_885 == 5'h15; // @[package.scala 31:81]
  assign _T_792_bits = {{3'd0}, _T_787}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _T_927_bits = _T_926 ? _T_792_bits : _T_925_bits; // @[package.scala 31:71]
  assign _T_927_rd = _T_926 ? io_in[11:7] : _T_925_rd; // @[package.scala 31:71]
  assign _T_927_rs1 = _T_926 ? 5'h2 : _T_925_rs1; // @[package.scala 31:71]
  assign _T_927_rs2 = _T_926 ? io_in[6:2] : _T_925_rs2; // @[package.scala 31:71]
  assign _T_927_rs3 = _T_926 ? io_in[31:27] : _T_925_rs3; // @[package.scala 31:71]
  assign _T_928 = _T_885 == 5'h16; // @[package.scala 31:81]
  assign _T_813_bits = {{4'd0}, _T_808}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _T_929_bits = _T_928 ? _T_813_bits : _T_927_bits; // @[package.scala 31:71]
  assign _T_929_rd = _T_928 ? io_in[11:7] : _T_927_rd; // @[package.scala 31:71]
  assign _T_929_rs1 = _T_928 ? 5'h2 : _T_927_rs1; // @[package.scala 31:71]
  assign _T_929_rs2 = _T_928 ? io_in[6:2] : _T_927_rs2; // @[package.scala 31:71]
  assign _T_929_rs3 = _T_928 ? io_in[31:27] : _T_927_rs3; // @[package.scala 31:71]
  assign _T_930 = _T_885 == 5'h17; // @[package.scala 31:81]
  assign _T_834_bits = {{3'd0}, _T_829}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _T_931_bits = _T_930 ? _T_834_bits : _T_929_bits; // @[package.scala 31:71]
  assign _T_931_rd = _T_930 ? io_in[11:7] : _T_929_rd; // @[package.scala 31:71]
  assign _T_931_rs1 = _T_930 ? 5'h2 : _T_929_rs1; // @[package.scala 31:71]
  assign _T_931_rs2 = _T_930 ? io_in[6:2] : _T_929_rs2; // @[package.scala 31:71]
  assign _T_931_rs3 = _T_930 ? io_in[31:27] : _T_929_rs3; // @[package.scala 31:71]
  assign _T_932 = _T_885 == 5'h18; // @[package.scala 31:81]
  assign _T_933_bits = _T_932 ? io_in : _T_931_bits; // @[package.scala 31:71]
  assign _T_933_rd = _T_932 ? io_in[11:7] : _T_931_rd; // @[package.scala 31:71]
  assign _T_933_rs1 = _T_932 ? io_in[19:15] : _T_931_rs1; // @[package.scala 31:71]
  assign _T_933_rs2 = _T_932 ? io_in[24:20] : _T_931_rs2; // @[package.scala 31:71]
  assign _T_933_rs3 = _T_932 ? io_in[31:27] : _T_931_rs3; // @[package.scala 31:71]
  assign _T_934 = _T_885 == 5'h19; // @[package.scala 31:81]
  assign _T_935_bits = _T_934 ? io_in : _T_933_bits; // @[package.scala 31:71]
  assign _T_935_rd = _T_934 ? io_in[11:7] : _T_933_rd; // @[package.scala 31:71]
  assign _T_935_rs1 = _T_934 ? io_in[19:15] : _T_933_rs1; // @[package.scala 31:71]
  assign _T_935_rs2 = _T_934 ? io_in[24:20] : _T_933_rs2; // @[package.scala 31:71]
  assign _T_935_rs3 = _T_934 ? io_in[31:27] : _T_933_rs3; // @[package.scala 31:71]
  assign _T_936 = _T_885 == 5'h1a; // @[package.scala 31:81]
  assign _T_937_bits = _T_936 ? io_in : _T_935_bits; // @[package.scala 31:71]
  assign _T_937_rd = _T_936 ? io_in[11:7] : _T_935_rd; // @[package.scala 31:71]
  assign _T_937_rs1 = _T_936 ? io_in[19:15] : _T_935_rs1; // @[package.scala 31:71]
  assign _T_937_rs2 = _T_936 ? io_in[24:20] : _T_935_rs2; // @[package.scala 31:71]
  assign _T_937_rs3 = _T_936 ? io_in[31:27] : _T_935_rs3; // @[package.scala 31:71]
  assign _T_938 = _T_885 == 5'h1b; // @[package.scala 31:81]
  assign _T_939_bits = _T_938 ? io_in : _T_937_bits; // @[package.scala 31:71]
  assign _T_939_rd = _T_938 ? io_in[11:7] : _T_937_rd; // @[package.scala 31:71]
  assign _T_939_rs1 = _T_938 ? io_in[19:15] : _T_937_rs1; // @[package.scala 31:71]
  assign _T_939_rs2 = _T_938 ? io_in[24:20] : _T_937_rs2; // @[package.scala 31:71]
  assign _T_939_rs3 = _T_938 ? io_in[31:27] : _T_937_rs3; // @[package.scala 31:71]
  assign _T_940 = _T_885 == 5'h1c; // @[package.scala 31:81]
  assign _T_941_bits = _T_940 ? io_in : _T_939_bits; // @[package.scala 31:71]
  assign _T_941_rd = _T_940 ? io_in[11:7] : _T_939_rd; // @[package.scala 31:71]
  assign _T_941_rs1 = _T_940 ? io_in[19:15] : _T_939_rs1; // @[package.scala 31:71]
  assign _T_941_rs2 = _T_940 ? io_in[24:20] : _T_939_rs2; // @[package.scala 31:71]
  assign _T_941_rs3 = _T_940 ? io_in[31:27] : _T_939_rs3; // @[package.scala 31:71]
  assign _T_942 = _T_885 == 5'h1d; // @[package.scala 31:81]
  assign _T_943_bits = _T_942 ? io_in : _T_941_bits; // @[package.scala 31:71]
  assign _T_943_rd = _T_942 ? io_in[11:7] : _T_941_rd; // @[package.scala 31:71]
  assign _T_943_rs1 = _T_942 ? io_in[19:15] : _T_941_rs1; // @[package.scala 31:71]
  assign _T_943_rs2 = _T_942 ? io_in[24:20] : _T_941_rs2; // @[package.scala 31:71]
  assign _T_943_rs3 = _T_942 ? io_in[31:27] : _T_941_rs3; // @[package.scala 31:71]
  assign _T_944 = _T_885 == 5'h1e; // @[package.scala 31:81]
  assign _T_945_bits = _T_944 ? io_in : _T_943_bits; // @[package.scala 31:71]
  assign _T_945_rd = _T_944 ? io_in[11:7] : _T_943_rd; // @[package.scala 31:71]
  assign _T_945_rs1 = _T_944 ? io_in[19:15] : _T_943_rs1; // @[package.scala 31:71]
  assign _T_945_rs2 = _T_944 ? io_in[24:20] : _T_943_rs2; // @[package.scala 31:71]
  assign _T_945_rs3 = _T_944 ? io_in[31:27] : _T_943_rs3; // @[package.scala 31:71]
  assign _T_946 = _T_885 == 5'h1f; // @[package.scala 31:81]
  assign io_out_bits = _T_946 ? io_in : _T_945_bits; // @[RVC.scala 164:12]
  assign io_out_rd = _T_946 ? io_in[11:7] : _T_945_rd; // @[RVC.scala 164:12]
  assign io_out_rs1 = _T_946 ? io_in[19:15] : _T_945_rs1; // @[RVC.scala 164:12]
  assign io_out_rs2 = _T_946 ? io_in[24:20] : _T_945_rs2; // @[RVC.scala 164:12]
  assign io_out_rs3 = _T_946 ? io_in[31:27] : _T_945_rs3; // @[RVC.scala 164:12]
  assign io_rvc = io_in[1:0] != 2'h3; // @[RVC.scala 163:12]
  assign RVCExpander_covSum = 30'h0;
  assign io_covSum = RVCExpander_covSum;
  assign metaAssert = 1'h0;
endmodule
module MulAddRecFNToRaw_preMul(
  input  [1:0]  io_op,
  input  [32:0] io_a,
  input  [32:0] io_b,
  input  [32:0] io_c,
  output [23:0] io_mulAddA,
  output [23:0] io_mulAddB,
  output [47:0] io_mulAddC,
  output        io_toPostMul_isSigNaNAny,
  output        io_toPostMul_isNaNAOrB,
  output        io_toPostMul_isInfA,
  output        io_toPostMul_isZeroA,
  output        io_toPostMul_isInfB,
  output        io_toPostMul_isZeroB,
  output        io_toPostMul_signProd,
  output        io_toPostMul_isNaNC,
  output        io_toPostMul_isInfC,
  output        io_toPostMul_isZeroC,
  output [9:0]  io_toPostMul_sExpSum,
  output        io_toPostMul_doSubMags,
  output        io_toPostMul_CIsDominant,
  output [4:0]  io_toPostMul_CDom_CAlignDist,
  output [25:0] io_toPostMul_highAlignedSigC,
  output        io_toPostMul_bit0AlignedSigC,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  rawA_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_16; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawA_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawA_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [24:0] rawA_sig; // @[Cat.scala 30:58]
  wire  rawB_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_33; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawB_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawB_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [24:0] rawB_sig; // @[Cat.scala 30:58]
  wire  rawC_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_50; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawC_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawC_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawC_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [24:0] rawC_sig; // @[Cat.scala 30:58]
  wire  _T_63; // @[MulAddRecFN.scala 98:30]
  wire  signProd; // @[MulAddRecFN.scala 98:42]
  wire [10:0] _T_65; // @[MulAddRecFN.scala 101:19]
  wire [10:0] sExpAlignedProd; // @[MulAddRecFN.scala 101:32]
  wire  _T_68; // @[MulAddRecFN.scala 103:30]
  wire  doSubMags; // @[MulAddRecFN.scala 103:42]
  wire [10:0] _GEN_0; // @[MulAddRecFN.scala 107:42]
  wire [10:0] sNatCAlignDist; // @[MulAddRecFN.scala 107:42]
  wire [9:0] posNatCAlignDist; // @[MulAddRecFN.scala 108:42]
  wire  _T_72; // @[MulAddRecFN.scala 109:35]
  wire  _T_73; // @[MulAddRecFN.scala 109:69]
  wire  isMinCAlign; // @[MulAddRecFN.scala 109:50]
  wire  _T_75; // @[MulAddRecFN.scala 111:60]
  wire  _T_76; // @[MulAddRecFN.scala 111:39]
  wire  CIsDominant; // @[MulAddRecFN.scala 111:23]
  wire  _T_77; // @[MulAddRecFN.scala 115:34]
  wire [6:0] _T_79; // @[MulAddRecFN.scala 115:16]
  wire [6:0] CAlignDist; // @[MulAddRecFN.scala 113:12]
  wire [24:0] _T_81; // @[MulAddRecFN.scala 121:16]
  wire [52:0] _T_83; // @[Bitwise.scala 72:12]
  wire [77:0] _T_85; // @[MulAddRecFN.scala 123:11]
  wire [77:0] mainAlignedSigC; // @[MulAddRecFN.scala 123:17]
  wire [26:0] _T_86; // @[MulAddRecFN.scala 125:30]
  wire  _T_101; // @[primitives.scala 121:54]
  wire  _T_103; // @[primitives.scala 121:54]
  wire  _T_105; // @[primitives.scala 121:54]
  wire  _T_107; // @[primitives.scala 121:54]
  wire  _T_109; // @[primitives.scala 121:54]
  wire  _T_111; // @[primitives.scala 121:54]
  wire  _T_113; // @[primitives.scala 124:57]
  wire [6:0] _T_119; // @[primitives.scala 125:20]
  wire [32:0] _T_121; // @[primitives.scala 77:58]
  wire [5:0] _T_137; // @[Cat.scala 30:58]
  wire [6:0] _GEN_1; // @[MulAddRecFN.scala 125:68]
  wire [6:0] _T_138; // @[MulAddRecFN.scala 125:68]
  wire  reduced4CExtra; // @[MulAddRecFN.scala 133:11]
  wire  _T_142; // @[MulAddRecFN.scala 137:39]
  wire  _T_144; // @[MulAddRecFN.scala 137:44]
  wire  _T_146; // @[MulAddRecFN.scala 138:39]
  wire  _T_147; // @[MulAddRecFN.scala 138:44]
  wire  _T_148; // @[MulAddRecFN.scala 136:16]
  wire [74:0] _T_149; // @[Cat.scala 30:58]
  wire [75:0] alignedSigC; // @[Cat.scala 30:58]
  wire  _T_153; // @[common.scala 81:46]
  wire  _T_156; // @[common.scala 81:46]
  wire  _T_157; // @[MulAddRecFN.scala 149:32]
  wire  _T_160; // @[common.scala 81:46]
  wire [10:0] _T_165; // @[MulAddRecFN.scala 161:53]
  wire [10:0] _T_166; // @[MulAddRecFN.scala 161:12]
  wire [29:0] MulAddRecFNToRaw_preMul_covSum;
  assign rawA_isZero = io_a[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_16 = io_a[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawA_isNaN = _T_16 & io_a[29]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawA_sign = io_a[32]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawA_sExp = {1'b0,$signed(io_a[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawA_sig = {1'h0,~rawA_isZero,io_a[22:0]}; // @[Cat.scala 30:58]
  assign rawB_isZero = io_b[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_33 = io_b[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawB_isNaN = _T_33 & io_b[29]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawB_sign = io_b[32]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawB_sExp = {1'b0,$signed(io_b[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawB_sig = {1'h0,~rawB_isZero,io_b[22:0]}; // @[Cat.scala 30:58]
  assign rawC_isZero = io_c[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_50 = io_c[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawC_isNaN = _T_50 & io_c[29]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawC_sign = io_c[32]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawC_sExp = {1'b0,$signed(io_c[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawC_sig = {1'h0,~rawC_isZero,io_c[22:0]}; // @[Cat.scala 30:58]
  assign _T_63 = rawA_sign ^ rawB_sign; // @[MulAddRecFN.scala 98:30]
  assign signProd = _T_63 ^ io_op[1]; // @[MulAddRecFN.scala 98:42]
  assign _T_65 = $signed(rawA_sExp) + $signed(rawB_sExp); // @[MulAddRecFN.scala 101:19]
  assign sExpAlignedProd = $signed(_T_65) + -11'she5; // @[MulAddRecFN.scala 101:32]
  assign _T_68 = signProd ^ rawC_sign; // @[MulAddRecFN.scala 103:30]
  assign doSubMags = _T_68 ^ io_op[0]; // @[MulAddRecFN.scala 103:42]
  assign _GEN_0 = {{1{rawC_sExp[9]}},rawC_sExp}; // @[MulAddRecFN.scala 107:42]
  assign sNatCAlignDist = $signed(sExpAlignedProd) - $signed(_GEN_0); // @[MulAddRecFN.scala 107:42]
  assign posNatCAlignDist = sNatCAlignDist[9:0]; // @[MulAddRecFN.scala 108:42]
  assign _T_72 = rawA_isZero | rawB_isZero; // @[MulAddRecFN.scala 109:35]
  assign _T_73 = $signed(sNatCAlignDist) < 11'sh0; // @[MulAddRecFN.scala 109:69]
  assign isMinCAlign = _T_72 | _T_73; // @[MulAddRecFN.scala 109:50]
  assign _T_75 = posNatCAlignDist <= 10'h18; // @[MulAddRecFN.scala 111:60]
  assign _T_76 = isMinCAlign | _T_75; // @[MulAddRecFN.scala 111:39]
  assign CIsDominant = ~rawC_isZero & _T_76; // @[MulAddRecFN.scala 111:23]
  assign _T_77 = posNatCAlignDist < 10'h4a; // @[MulAddRecFN.scala 115:34]
  assign _T_79 = _T_77 ? posNatCAlignDist[6:0] : 7'h4a; // @[MulAddRecFN.scala 115:16]
  assign CAlignDist = isMinCAlign ? 7'h0 : _T_79; // @[MulAddRecFN.scala 113:12]
  assign _T_81 = doSubMags ? ~rawC_sig : rawC_sig; // @[MulAddRecFN.scala 121:16]
  assign _T_83 = doSubMags ? 53'h1fffffffffffff : 53'h0; // @[Bitwise.scala 72:12]
  assign _T_85 = {_T_81,_T_83}; // @[MulAddRecFN.scala 123:11]
  assign mainAlignedSigC = $signed(_T_85) >>> CAlignDist; // @[MulAddRecFN.scala 123:17]
  assign _T_86 = {rawC_sig, 2'h0}; // @[MulAddRecFN.scala 125:30]
  assign _T_101 = _T_86[3:0] != 4'h0; // @[primitives.scala 121:54]
  assign _T_103 = _T_86[7:4] != 4'h0; // @[primitives.scala 121:54]
  assign _T_105 = _T_86[11:8] != 4'h0; // @[primitives.scala 121:54]
  assign _T_107 = _T_86[15:12] != 4'h0; // @[primitives.scala 121:54]
  assign _T_109 = _T_86[19:16] != 4'h0; // @[primitives.scala 121:54]
  assign _T_111 = _T_86[23:20] != 4'h0; // @[primitives.scala 121:54]
  assign _T_113 = _T_86[26:24] != 3'h0; // @[primitives.scala 124:57]
  assign _T_119 = {_T_113,_T_111,_T_109,_T_107,_T_105,_T_103,_T_101}; // @[primitives.scala 125:20]
  assign _T_121 = -33'sh100000000 >>> CAlignDist[6:2]; // @[primitives.scala 77:58]
  assign _T_137 = {_T_121[14],_T_121[15],_T_121[16],_T_121[17],_T_121[18],_T_121[19]}; // @[Cat.scala 30:58]
  assign _GEN_1 = {{1'd0}, _T_137}; // @[MulAddRecFN.scala 125:68]
  assign _T_138 = _T_119 & _GEN_1; // @[MulAddRecFN.scala 125:68]
  assign reduced4CExtra = _T_138 != 7'h0; // @[MulAddRecFN.scala 133:11]
  assign _T_142 = ~mainAlignedSigC[2:0] == 3'h0; // @[MulAddRecFN.scala 137:39]
  assign _T_144 = _T_142 & ~reduced4CExtra; // @[MulAddRecFN.scala 137:44]
  assign _T_146 = mainAlignedSigC[2:0] != 3'h0; // @[MulAddRecFN.scala 138:39]
  assign _T_147 = _T_146 | reduced4CExtra; // @[MulAddRecFN.scala 138:44]
  assign _T_148 = doSubMags ? _T_144 : _T_147; // @[MulAddRecFN.scala 136:16]
  assign _T_149 = mainAlignedSigC[77:3]; // @[Cat.scala 30:58]
  assign alignedSigC = {_T_149,_T_148}; // @[Cat.scala 30:58]
  assign _T_153 = rawA_isNaN & ~rawA_sig[22]; // @[common.scala 81:46]
  assign _T_156 = rawB_isNaN & ~rawB_sig[22]; // @[common.scala 81:46]
  assign _T_157 = _T_153 | _T_156; // @[MulAddRecFN.scala 149:32]
  assign _T_160 = rawC_isNaN & ~rawC_sig[22]; // @[common.scala 81:46]
  assign _T_165 = $signed(sExpAlignedProd) - 11'sh18; // @[MulAddRecFN.scala 161:53]
  assign _T_166 = CIsDominant ? $signed({{1{rawC_sExp[9]}},rawC_sExp}) : $signed(_T_165); // @[MulAddRecFN.scala 161:12]
  assign io_mulAddA = rawA_sig[23:0]; // @[MulAddRecFN.scala 144:16]
  assign io_mulAddB = rawB_sig[23:0]; // @[MulAddRecFN.scala 145:16]
  assign io_mulAddC = alignedSigC[48:1]; // @[MulAddRecFN.scala 146:16]
  assign io_toPostMul_isSigNaNAny = _T_157 | _T_160; // @[MulAddRecFN.scala 148:30]
  assign io_toPostMul_isNaNAOrB = rawA_isNaN | rawB_isNaN; // @[MulAddRecFN.scala 151:28]
  assign io_toPostMul_isInfA = _T_16 & ~io_a[29]; // @[MulAddRecFN.scala 152:28]
  assign io_toPostMul_isZeroA = io_a[31:29] == 3'h0; // @[MulAddRecFN.scala 153:28]
  assign io_toPostMul_isInfB = _T_33 & ~io_b[29]; // @[MulAddRecFN.scala 154:28]
  assign io_toPostMul_isZeroB = io_b[31:29] == 3'h0; // @[MulAddRecFN.scala 155:28]
  assign io_toPostMul_signProd = _T_63 ^ io_op[1]; // @[MulAddRecFN.scala 156:28]
  assign io_toPostMul_isNaNC = _T_50 & io_c[29]; // @[MulAddRecFN.scala 157:28]
  assign io_toPostMul_isInfC = _T_50 & ~io_c[29]; // @[MulAddRecFN.scala 158:28]
  assign io_toPostMul_isZeroC = io_c[31:29] == 3'h0; // @[MulAddRecFN.scala 159:28]
  assign io_toPostMul_sExpSum = _T_166[9:0]; // @[MulAddRecFN.scala 160:28]
  assign io_toPostMul_doSubMags = _T_68 ^ io_op[0]; // @[MulAddRecFN.scala 162:28]
  assign io_toPostMul_CIsDominant = ~rawC_isZero & _T_76; // @[MulAddRecFN.scala 163:30]
  assign io_toPostMul_CDom_CAlignDist = CAlignDist[4:0]; // @[MulAddRecFN.scala 164:34]
  assign io_toPostMul_highAlignedSigC = alignedSigC[74:49]; // @[MulAddRecFN.scala 165:34]
  assign io_toPostMul_bit0AlignedSigC = alignedSigC[0]; // @[MulAddRecFN.scala 167:34]
  assign MulAddRecFNToRaw_preMul_covSum = 30'h0;
  assign io_covSum = MulAddRecFNToRaw_preMul_covSum;
  assign metaAssert = 1'h0;
endmodule
module MulAddRecFNToRaw_postMul(
  input         io_fromPreMul_isSigNaNAny,
  input         io_fromPreMul_isNaNAOrB,
  input         io_fromPreMul_isInfA,
  input         io_fromPreMul_isZeroA,
  input         io_fromPreMul_isInfB,
  input         io_fromPreMul_isZeroB,
  input         io_fromPreMul_signProd,
  input         io_fromPreMul_isNaNC,
  input         io_fromPreMul_isInfC,
  input         io_fromPreMul_isZeroC,
  input  [9:0]  io_fromPreMul_sExpSum,
  input         io_fromPreMul_doSubMags,
  input         io_fromPreMul_CIsDominant,
  input  [4:0]  io_fromPreMul_CDom_CAlignDist,
  input  [25:0] io_fromPreMul_highAlignedSigC,
  input         io_fromPreMul_bit0AlignedSigC,
  input  [48:0] io_mulAddResult,
  input  [2:0]  io_roundingMode,
  output        io_invalidExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [9:0]  io_rawOut_sExp,
  output [26:0] io_rawOut_sig,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundingMode_min; // @[MulAddRecFN.scala 188:45]
  wire  CDom_sign; // @[MulAddRecFN.scala 192:42]
  wire [25:0] _T_11; // @[MulAddRecFN.scala 195:47]
  wire [25:0] _T_12; // @[MulAddRecFN.scala 194:16]
  wire [74:0] sigSum; // @[Cat.scala 30:58]
  wire [1:0] _T_15; // @[MulAddRecFN.scala 205:69]
  wire [9:0] _GEN_0; // @[MulAddRecFN.scala 205:43]
  wire [9:0] CDom_sExp; // @[MulAddRecFN.scala 205:43]
  wire [49:0] _T_23; // @[Cat.scala 30:58]
  wire [49:0] CDom_absSigSum; // @[MulAddRecFN.scala 207:12]
  wire  _T_26; // @[MulAddRecFN.scala 217:36]
  wire  _T_28; // @[MulAddRecFN.scala 218:37]
  wire  CDom_absSigSumExtra; // @[MulAddRecFN.scala 216:12]
  wire [80:0] _GEN_1; // @[MulAddRecFN.scala 221:24]
  wire [80:0] _T_29; // @[MulAddRecFN.scala 221:24]
  wire [28:0] CDom_mainSig; // @[MulAddRecFN.scala 221:56]
  wire [26:0] _T_31; // @[MulAddRecFN.scala 224:53]
  wire  _T_46; // @[primitives.scala 121:54]
  wire  _T_48; // @[primitives.scala 121:54]
  wire  _T_50; // @[primitives.scala 121:54]
  wire  _T_52; // @[primitives.scala 121:54]
  wire  _T_54; // @[primitives.scala 121:54]
  wire  _T_56; // @[primitives.scala 121:54]
  wire  _T_58; // @[primitives.scala 124:57]
  wire [6:0] _T_64; // @[primitives.scala 125:20]
  wire [8:0] _T_67; // @[primitives.scala 77:58]
  wire [5:0] _T_83; // @[Cat.scala 30:58]
  wire [6:0] _GEN_2; // @[MulAddRecFN.scala 224:72]
  wire [6:0] _T_84; // @[MulAddRecFN.scala 224:72]
  wire  CDom_reduced4SigExtra; // @[MulAddRecFN.scala 225:73]
  wire  _T_87; // @[MulAddRecFN.scala 228:32]
  wire  _T_88; // @[MulAddRecFN.scala 228:36]
  wire  _T_89; // @[MulAddRecFN.scala 228:61]
  wire [26:0] CDom_sig; // @[Cat.scala 30:58]
  wire  notCDom_signSigSum; // @[MulAddRecFN.scala 234:36]
  wire [50:0] _GEN_3; // @[MulAddRecFN.scala 238:41]
  wire [50:0] _T_94; // @[MulAddRecFN.scala 238:41]
  wire [50:0] notCDom_absSigSum; // @[MulAddRecFN.scala 236:12]
  wire  _T_128; // @[primitives.scala 104:54]
  wire  _T_130; // @[primitives.scala 104:54]
  wire  _T_132; // @[primitives.scala 104:54]
  wire  _T_134; // @[primitives.scala 104:54]
  wire  _T_136; // @[primitives.scala 104:54]
  wire  _T_138; // @[primitives.scala 104:54]
  wire  _T_140; // @[primitives.scala 104:54]
  wire  _T_142; // @[primitives.scala 104:54]
  wire  _T_144; // @[primitives.scala 104:54]
  wire  _T_146; // @[primitives.scala 104:54]
  wire  _T_148; // @[primitives.scala 104:54]
  wire  _T_150; // @[primitives.scala 104:54]
  wire  _T_152; // @[primitives.scala 104:54]
  wire  _T_154; // @[primitives.scala 104:54]
  wire  _T_156; // @[primitives.scala 104:54]
  wire  _T_158; // @[primitives.scala 104:54]
  wire  _T_160; // @[primitives.scala 104:54]
  wire  _T_162; // @[primitives.scala 104:54]
  wire  _T_164; // @[primitives.scala 104:54]
  wire  _T_166; // @[primitives.scala 104:54]
  wire  _T_168; // @[primitives.scala 104:54]
  wire  _T_170; // @[primitives.scala 104:54]
  wire  _T_172; // @[primitives.scala 104:54]
  wire  _T_174; // @[primitives.scala 104:54]
  wire  _T_176; // @[primitives.scala 104:54]
  wire [5:0] _T_183; // @[primitives.scala 108:20]
  wire [12:0] _T_190; // @[primitives.scala 108:20]
  wire [5:0] _T_195; // @[primitives.scala 108:20]
  wire [25:0] notCDom_reduced2AbsSigSum; // @[primitives.scala 108:20]
  wire [15:0] _T_207; // @[Bitwise.scala 103:31]
  wire [15:0] _T_209; // @[Bitwise.scala 103:65]
  wire [15:0] _T_211; // @[Bitwise.scala 103:75]
  wire [15:0] _T_212; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_4; // @[Bitwise.scala 103:31]
  wire [15:0] _T_217; // @[Bitwise.scala 103:31]
  wire [15:0] _T_219; // @[Bitwise.scala 103:65]
  wire [15:0] _T_221; // @[Bitwise.scala 103:75]
  wire [15:0] _T_222; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_5; // @[Bitwise.scala 103:31]
  wire [15:0] _T_227; // @[Bitwise.scala 103:31]
  wire [15:0] _T_229; // @[Bitwise.scala 103:65]
  wire [15:0] _T_231; // @[Bitwise.scala 103:75]
  wire [15:0] _T_232; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_6; // @[Bitwise.scala 103:31]
  wire [15:0] _T_237; // @[Bitwise.scala 103:31]
  wire [15:0] _T_239; // @[Bitwise.scala 103:65]
  wire [15:0] _T_241; // @[Bitwise.scala 103:75]
  wire [15:0] _T_242; // @[Bitwise.scala 103:39]
  wire [7:0] _T_248; // @[Bitwise.scala 103:31]
  wire [7:0] _T_250; // @[Bitwise.scala 103:65]
  wire [7:0] _T_252; // @[Bitwise.scala 103:75]
  wire [7:0] _T_253; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_7; // @[Bitwise.scala 103:31]
  wire [7:0] _T_258; // @[Bitwise.scala 103:31]
  wire [7:0] _T_260; // @[Bitwise.scala 103:65]
  wire [7:0] _T_262; // @[Bitwise.scala 103:75]
  wire [7:0] _T_263; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_8; // @[Bitwise.scala 103:31]
  wire [7:0] _T_268; // @[Bitwise.scala 103:31]
  wire [7:0] _T_270; // @[Bitwise.scala 103:65]
  wire [7:0] _T_272; // @[Bitwise.scala 103:75]
  wire [7:0] _T_273; // @[Bitwise.scala 103:39]
  wire [25:0] _T_279; // @[Cat.scala 30:58]
  wire [4:0] _T_306; // @[Mux.scala 31:69]
  wire [4:0] _T_307; // @[Mux.scala 31:69]
  wire [4:0] _T_308; // @[Mux.scala 31:69]
  wire [4:0] _T_309; // @[Mux.scala 31:69]
  wire [4:0] _T_310; // @[Mux.scala 31:69]
  wire [4:0] _T_311; // @[Mux.scala 31:69]
  wire [4:0] _T_312; // @[Mux.scala 31:69]
  wire [4:0] _T_313; // @[Mux.scala 31:69]
  wire [4:0] _T_314; // @[Mux.scala 31:69]
  wire [4:0] _T_315; // @[Mux.scala 31:69]
  wire [4:0] _T_316; // @[Mux.scala 31:69]
  wire [4:0] _T_317; // @[Mux.scala 31:69]
  wire [4:0] _T_318; // @[Mux.scala 31:69]
  wire [4:0] _T_319; // @[Mux.scala 31:69]
  wire [4:0] _T_320; // @[Mux.scala 31:69]
  wire [4:0] _T_321; // @[Mux.scala 31:69]
  wire [4:0] _T_322; // @[Mux.scala 31:69]
  wire [4:0] _T_323; // @[Mux.scala 31:69]
  wire [4:0] _T_324; // @[Mux.scala 31:69]
  wire [4:0] _T_325; // @[Mux.scala 31:69]
  wire [4:0] _T_326; // @[Mux.scala 31:69]
  wire [4:0] _T_327; // @[Mux.scala 31:69]
  wire [4:0] _T_328; // @[Mux.scala 31:69]
  wire [4:0] _T_329; // @[Mux.scala 31:69]
  wire [4:0] notCDom_normDistReduced2; // @[Mux.scala 31:69]
  wire [5:0] notCDom_nearNormDist; // @[MulAddRecFN.scala 242:56]
  wire [6:0] _T_330; // @[MulAddRecFN.scala 243:69]
  wire [9:0] _GEN_9; // @[MulAddRecFN.scala 243:46]
  wire [9:0] notCDom_sExp; // @[MulAddRecFN.scala 243:46]
  wire [113:0] _GEN_10; // @[MulAddRecFN.scala 245:27]
  wire [113:0] _T_333; // @[MulAddRecFN.scala 245:27]
  wire [28:0] notCDom_mainSig; // @[MulAddRecFN.scala 245:50]
  wire  _T_350; // @[primitives.scala 104:54]
  wire  _T_352; // @[primitives.scala 104:54]
  wire  _T_354; // @[primitives.scala 104:54]
  wire  _T_356; // @[primitives.scala 104:54]
  wire  _T_358; // @[primitives.scala 104:54]
  wire  _T_360; // @[primitives.scala 104:54]
  wire [6:0] _T_368; // @[primitives.scala 108:20]
  wire [16:0] _T_371; // @[primitives.scala 77:58]
  wire [5:0] _T_387; // @[Cat.scala 30:58]
  wire [6:0] _GEN_11; // @[MulAddRecFN.scala 249:78]
  wire [6:0] _T_388; // @[MulAddRecFN.scala 249:78]
  wire  notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 251:11]
  wire  _T_391; // @[MulAddRecFN.scala 254:35]
  wire  _T_392; // @[MulAddRecFN.scala 254:39]
  wire [26:0] notCDom_sig; // @[Cat.scala 30:58]
  wire  notCDom_completeCancellation; // @[MulAddRecFN.scala 257:50]
  wire  _T_394; // @[MulAddRecFN.scala 261:36]
  wire  notCDom_sign; // @[MulAddRecFN.scala 259:12]
  wire  notNaN_isInfProd; // @[MulAddRecFN.scala 266:49]
  wire  notNaN_isInfOut; // @[MulAddRecFN.scala 267:44]
  wire  _T_395; // @[MulAddRecFN.scala 269:32]
  wire  notNaN_addZeros; // @[MulAddRecFN.scala 269:58]
  wire  _T_396; // @[MulAddRecFN.scala 274:31]
  wire  _T_397; // @[MulAddRecFN.scala 273:35]
  wire  _T_398; // @[MulAddRecFN.scala 275:32]
  wire  _T_399; // @[MulAddRecFN.scala 274:57]
  wire  _T_402; // @[MulAddRecFN.scala 276:36]
  wire  _T_403; // @[MulAddRecFN.scala 277:61]
  wire  _T_404; // @[MulAddRecFN.scala 278:35]
  wire  _T_408; // @[MulAddRecFN.scala 285:42]
  wire  _T_410; // @[MulAddRecFN.scala 287:27]
  wire  _T_411; // @[MulAddRecFN.scala 288:31]
  wire  _T_412; // @[MulAddRecFN.scala 287:54]
  wire  _T_414; // @[MulAddRecFN.scala 289:26]
  wire  _T_415; // @[MulAddRecFN.scala 289:48]
  wire  _T_416; // @[MulAddRecFN.scala 290:36]
  wire  _T_417; // @[MulAddRecFN.scala 288:43]
  wire  _T_418; // @[MulAddRecFN.scala 291:26]
  wire  _T_419; // @[MulAddRecFN.scala 292:37]
  wire  _T_420; // @[MulAddRecFN.scala 291:46]
  wire  _T_421; // @[MulAddRecFN.scala 290:48]
  wire  _T_424; // @[MulAddRecFN.scala 293:28]
  wire  _T_425; // @[MulAddRecFN.scala 294:17]
  wire  _T_426; // @[MulAddRecFN.scala 293:49]
  wire [29:0] MulAddRecFNToRaw_postMul_covSum;
  assign roundingMode_min = io_roundingMode == 3'h2; // @[MulAddRecFN.scala 188:45]
  assign CDom_sign = io_fromPreMul_signProd ^ io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 192:42]
  assign _T_11 = io_fromPreMul_highAlignedSigC + 26'h1; // @[MulAddRecFN.scala 195:47]
  assign _T_12 = io_mulAddResult[48] ? _T_11 : io_fromPreMul_highAlignedSigC; // @[MulAddRecFN.scala 194:16]
  assign sigSum = {_T_12,io_mulAddResult[47:0],io_fromPreMul_bit0AlignedSigC}; // @[Cat.scala 30:58]
  assign _T_15 = {1'b0,$signed(io_fromPreMul_doSubMags)}; // @[MulAddRecFN.scala 205:69]
  assign _GEN_0 = {{8{_T_15[1]}},_T_15}; // @[MulAddRecFN.scala 205:43]
  assign CDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_0); // @[MulAddRecFN.scala 205:43]
  assign _T_23 = {1'h0,io_fromPreMul_highAlignedSigC[25:24],sigSum[72:26]}; // @[Cat.scala 30:58]
  assign CDom_absSigSum = io_fromPreMul_doSubMags ? ~sigSum[74:25] : _T_23; // @[MulAddRecFN.scala 207:12]
  assign _T_26 = ~sigSum[24:1] != 24'h0; // @[MulAddRecFN.scala 217:36]
  assign _T_28 = sigSum[25:1] != 25'h0; // @[MulAddRecFN.scala 218:37]
  assign CDom_absSigSumExtra = io_fromPreMul_doSubMags ? _T_26 : _T_28; // @[MulAddRecFN.scala 216:12]
  assign _GEN_1 = {{31'd0}, CDom_absSigSum}; // @[MulAddRecFN.scala 221:24]
  assign _T_29 = _GEN_1 << io_fromPreMul_CDom_CAlignDist; // @[MulAddRecFN.scala 221:24]
  assign CDom_mainSig = _T_29[49:21]; // @[MulAddRecFN.scala 221:56]
  assign _T_31 = {CDom_absSigSum[23:0], 3'h0}; // @[MulAddRecFN.scala 224:53]
  assign _T_46 = _T_31[3:0] != 4'h0; // @[primitives.scala 121:54]
  assign _T_48 = _T_31[7:4] != 4'h0; // @[primitives.scala 121:54]
  assign _T_50 = _T_31[11:8] != 4'h0; // @[primitives.scala 121:54]
  assign _T_52 = _T_31[15:12] != 4'h0; // @[primitives.scala 121:54]
  assign _T_54 = _T_31[19:16] != 4'h0; // @[primitives.scala 121:54]
  assign _T_56 = _T_31[23:20] != 4'h0; // @[primitives.scala 121:54]
  assign _T_58 = _T_31[26:24] != 3'h0; // @[primitives.scala 124:57]
  assign _T_64 = {_T_58,_T_56,_T_54,_T_52,_T_50,_T_48,_T_46}; // @[primitives.scala 125:20]
  assign _T_67 = -9'sh100 >>> ~io_fromPreMul_CDom_CAlignDist[4:2]; // @[primitives.scala 77:58]
  assign _T_83 = {_T_67[1],_T_67[2],_T_67[3],_T_67[4],_T_67[5],_T_67[6]}; // @[Cat.scala 30:58]
  assign _GEN_2 = {{1'd0}, _T_83}; // @[MulAddRecFN.scala 224:72]
  assign _T_84 = _T_64 & _GEN_2; // @[MulAddRecFN.scala 224:72]
  assign CDom_reduced4SigExtra = _T_84 != 7'h0; // @[MulAddRecFN.scala 225:73]
  assign _T_87 = CDom_mainSig[2:0] != 3'h0; // @[MulAddRecFN.scala 228:32]
  assign _T_88 = _T_87 | CDom_reduced4SigExtra; // @[MulAddRecFN.scala 228:36]
  assign _T_89 = _T_88 | CDom_absSigSumExtra; // @[MulAddRecFN.scala 228:61]
  assign CDom_sig = {CDom_mainSig[28:3],_T_89}; // @[Cat.scala 30:58]
  assign notCDom_signSigSum = sigSum[51]; // @[MulAddRecFN.scala 234:36]
  assign _GEN_3 = {{50'd0}, io_fromPreMul_doSubMags}; // @[MulAddRecFN.scala 238:41]
  assign _T_94 = sigSum[50:0] + _GEN_3; // @[MulAddRecFN.scala 238:41]
  assign notCDom_absSigSum = notCDom_signSigSum ? ~sigSum[50:0] : _T_94; // @[MulAddRecFN.scala 236:12]
  assign _T_128 = notCDom_absSigSum[1:0] != 2'h0; // @[primitives.scala 104:54]
  assign _T_130 = notCDom_absSigSum[3:2] != 2'h0; // @[primitives.scala 104:54]
  assign _T_132 = notCDom_absSigSum[5:4] != 2'h0; // @[primitives.scala 104:54]
  assign _T_134 = notCDom_absSigSum[7:6] != 2'h0; // @[primitives.scala 104:54]
  assign _T_136 = notCDom_absSigSum[9:8] != 2'h0; // @[primitives.scala 104:54]
  assign _T_138 = notCDom_absSigSum[11:10] != 2'h0; // @[primitives.scala 104:54]
  assign _T_140 = notCDom_absSigSum[13:12] != 2'h0; // @[primitives.scala 104:54]
  assign _T_142 = notCDom_absSigSum[15:14] != 2'h0; // @[primitives.scala 104:54]
  assign _T_144 = notCDom_absSigSum[17:16] != 2'h0; // @[primitives.scala 104:54]
  assign _T_146 = notCDom_absSigSum[19:18] != 2'h0; // @[primitives.scala 104:54]
  assign _T_148 = notCDom_absSigSum[21:20] != 2'h0; // @[primitives.scala 104:54]
  assign _T_150 = notCDom_absSigSum[23:22] != 2'h0; // @[primitives.scala 104:54]
  assign _T_152 = notCDom_absSigSum[25:24] != 2'h0; // @[primitives.scala 104:54]
  assign _T_154 = notCDom_absSigSum[27:26] != 2'h0; // @[primitives.scala 104:54]
  assign _T_156 = notCDom_absSigSum[29:28] != 2'h0; // @[primitives.scala 104:54]
  assign _T_158 = notCDom_absSigSum[31:30] != 2'h0; // @[primitives.scala 104:54]
  assign _T_160 = notCDom_absSigSum[33:32] != 2'h0; // @[primitives.scala 104:54]
  assign _T_162 = notCDom_absSigSum[35:34] != 2'h0; // @[primitives.scala 104:54]
  assign _T_164 = notCDom_absSigSum[37:36] != 2'h0; // @[primitives.scala 104:54]
  assign _T_166 = notCDom_absSigSum[39:38] != 2'h0; // @[primitives.scala 104:54]
  assign _T_168 = notCDom_absSigSum[41:40] != 2'h0; // @[primitives.scala 104:54]
  assign _T_170 = notCDom_absSigSum[43:42] != 2'h0; // @[primitives.scala 104:54]
  assign _T_172 = notCDom_absSigSum[45:44] != 2'h0; // @[primitives.scala 104:54]
  assign _T_174 = notCDom_absSigSum[47:46] != 2'h0; // @[primitives.scala 104:54]
  assign _T_176 = notCDom_absSigSum[49:48] != 2'h0; // @[primitives.scala 104:54]
  assign _T_183 = {_T_138,_T_136,_T_134,_T_132,_T_130,_T_128}; // @[primitives.scala 108:20]
  assign _T_190 = {_T_152,_T_150,_T_148,_T_146,_T_144,_T_142,_T_140,_T_183}; // @[primitives.scala 108:20]
  assign _T_195 = {_T_164,_T_162,_T_160,_T_158,_T_156,_T_154}; // @[primitives.scala 108:20]
  assign notCDom_reduced2AbsSigSum = {notCDom_absSigSum[50],_T_176,_T_174,_T_172,_T_170,_T_168,_T_166,_T_195,_T_190}; // @[primitives.scala 108:20]
  assign _T_207 = {{8'd0}, notCDom_reduced2AbsSigSum[15:8]}; // @[Bitwise.scala 103:31]
  assign _T_209 = {notCDom_reduced2AbsSigSum[7:0], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_211 = _T_209 & 16'hff00; // @[Bitwise.scala 103:75]
  assign _T_212 = _T_207 | _T_211; // @[Bitwise.scala 103:39]
  assign _GEN_4 = {{4'd0}, _T_212[15:4]}; // @[Bitwise.scala 103:31]
  assign _T_217 = _GEN_4 & 16'hf0f; // @[Bitwise.scala 103:31]
  assign _T_219 = {_T_212[11:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_221 = _T_219 & 16'hf0f0; // @[Bitwise.scala 103:75]
  assign _T_222 = _T_217 | _T_221; // @[Bitwise.scala 103:39]
  assign _GEN_5 = {{2'd0}, _T_222[15:2]}; // @[Bitwise.scala 103:31]
  assign _T_227 = _GEN_5 & 16'h3333; // @[Bitwise.scala 103:31]
  assign _T_229 = {_T_222[13:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_231 = _T_229 & 16'hcccc; // @[Bitwise.scala 103:75]
  assign _T_232 = _T_227 | _T_231; // @[Bitwise.scala 103:39]
  assign _GEN_6 = {{1'd0}, _T_232[15:1]}; // @[Bitwise.scala 103:31]
  assign _T_237 = _GEN_6 & 16'h5555; // @[Bitwise.scala 103:31]
  assign _T_239 = {_T_232[14:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_241 = _T_239 & 16'haaaa; // @[Bitwise.scala 103:75]
  assign _T_242 = _T_237 | _T_241; // @[Bitwise.scala 103:39]
  assign _T_248 = {{4'd0}, notCDom_reduced2AbsSigSum[23:20]}; // @[Bitwise.scala 103:31]
  assign _T_250 = {notCDom_reduced2AbsSigSum[19:16], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_252 = _T_250 & 8'hf0; // @[Bitwise.scala 103:75]
  assign _T_253 = _T_248 | _T_252; // @[Bitwise.scala 103:39]
  assign _GEN_7 = {{2'd0}, _T_253[7:2]}; // @[Bitwise.scala 103:31]
  assign _T_258 = _GEN_7 & 8'h33; // @[Bitwise.scala 103:31]
  assign _T_260 = {_T_253[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_262 = _T_260 & 8'hcc; // @[Bitwise.scala 103:75]
  assign _T_263 = _T_258 | _T_262; // @[Bitwise.scala 103:39]
  assign _GEN_8 = {{1'd0}, _T_263[7:1]}; // @[Bitwise.scala 103:31]
  assign _T_268 = _GEN_8 & 8'h55; // @[Bitwise.scala 103:31]
  assign _T_270 = {_T_263[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_272 = _T_270 & 8'haa; // @[Bitwise.scala 103:75]
  assign _T_273 = _T_268 | _T_272; // @[Bitwise.scala 103:39]
  assign _T_279 = {_T_242,_T_273,notCDom_reduced2AbsSigSum[24],notCDom_reduced2AbsSigSum[25]}; // @[Cat.scala 30:58]
  assign _T_306 = _T_279[24] ? 5'h18 : 5'h19; // @[Mux.scala 31:69]
  assign _T_307 = _T_279[23] ? 5'h17 : _T_306; // @[Mux.scala 31:69]
  assign _T_308 = _T_279[22] ? 5'h16 : _T_307; // @[Mux.scala 31:69]
  assign _T_309 = _T_279[21] ? 5'h15 : _T_308; // @[Mux.scala 31:69]
  assign _T_310 = _T_279[20] ? 5'h14 : _T_309; // @[Mux.scala 31:69]
  assign _T_311 = _T_279[19] ? 5'h13 : _T_310; // @[Mux.scala 31:69]
  assign _T_312 = _T_279[18] ? 5'h12 : _T_311; // @[Mux.scala 31:69]
  assign _T_313 = _T_279[17] ? 5'h11 : _T_312; // @[Mux.scala 31:69]
  assign _T_314 = _T_279[16] ? 5'h10 : _T_313; // @[Mux.scala 31:69]
  assign _T_315 = _T_279[15] ? 5'hf : _T_314; // @[Mux.scala 31:69]
  assign _T_316 = _T_279[14] ? 5'he : _T_315; // @[Mux.scala 31:69]
  assign _T_317 = _T_279[13] ? 5'hd : _T_316; // @[Mux.scala 31:69]
  assign _T_318 = _T_279[12] ? 5'hc : _T_317; // @[Mux.scala 31:69]
  assign _T_319 = _T_279[11] ? 5'hb : _T_318; // @[Mux.scala 31:69]
  assign _T_320 = _T_279[10] ? 5'ha : _T_319; // @[Mux.scala 31:69]
  assign _T_321 = _T_279[9] ? 5'h9 : _T_320; // @[Mux.scala 31:69]
  assign _T_322 = _T_279[8] ? 5'h8 : _T_321; // @[Mux.scala 31:69]
  assign _T_323 = _T_279[7] ? 5'h7 : _T_322; // @[Mux.scala 31:69]
  assign _T_324 = _T_279[6] ? 5'h6 : _T_323; // @[Mux.scala 31:69]
  assign _T_325 = _T_279[5] ? 5'h5 : _T_324; // @[Mux.scala 31:69]
  assign _T_326 = _T_279[4] ? 5'h4 : _T_325; // @[Mux.scala 31:69]
  assign _T_327 = _T_279[3] ? 5'h3 : _T_326; // @[Mux.scala 31:69]
  assign _T_328 = _T_279[2] ? 5'h2 : _T_327; // @[Mux.scala 31:69]
  assign _T_329 = _T_279[1] ? 5'h1 : _T_328; // @[Mux.scala 31:69]
  assign notCDom_normDistReduced2 = _T_279[0] ? 5'h0 : _T_329; // @[Mux.scala 31:69]
  assign notCDom_nearNormDist = {notCDom_normDistReduced2, 1'h0}; // @[MulAddRecFN.scala 242:56]
  assign _T_330 = {1'b0,$signed(notCDom_nearNormDist)}; // @[MulAddRecFN.scala 243:69]
  assign _GEN_9 = {{3{_T_330[6]}},_T_330}; // @[MulAddRecFN.scala 243:46]
  assign notCDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_9); // @[MulAddRecFN.scala 243:46]
  assign _GEN_10 = {{63'd0}, notCDom_absSigSum}; // @[MulAddRecFN.scala 245:27]
  assign _T_333 = _GEN_10 << notCDom_nearNormDist; // @[MulAddRecFN.scala 245:27]
  assign notCDom_mainSig = _T_333[51:23]; // @[MulAddRecFN.scala 245:50]
  assign _T_350 = notCDom_reduced2AbsSigSum[1:0] != 2'h0; // @[primitives.scala 104:54]
  assign _T_352 = notCDom_reduced2AbsSigSum[3:2] != 2'h0; // @[primitives.scala 104:54]
  assign _T_354 = notCDom_reduced2AbsSigSum[5:4] != 2'h0; // @[primitives.scala 104:54]
  assign _T_356 = notCDom_reduced2AbsSigSum[7:6] != 2'h0; // @[primitives.scala 104:54]
  assign _T_358 = notCDom_reduced2AbsSigSum[9:8] != 2'h0; // @[primitives.scala 104:54]
  assign _T_360 = notCDom_reduced2AbsSigSum[11:10] != 2'h0; // @[primitives.scala 104:54]
  assign _T_368 = {notCDom_reduced2AbsSigSum[12],_T_360,_T_358,_T_356,_T_354,_T_352,_T_350}; // @[primitives.scala 108:20]
  assign _T_371 = -17'sh10000 >>> ~notCDom_normDistReduced2[4:1]; // @[primitives.scala 77:58]
  assign _T_387 = {_T_371[1],_T_371[2],_T_371[3],_T_371[4],_T_371[5],_T_371[6]}; // @[Cat.scala 30:58]
  assign _GEN_11 = {{1'd0}, _T_387}; // @[MulAddRecFN.scala 249:78]
  assign _T_388 = _T_368 & _GEN_11; // @[MulAddRecFN.scala 249:78]
  assign notCDom_reduced4SigExtra = _T_388 != 7'h0; // @[MulAddRecFN.scala 251:11]
  assign _T_391 = notCDom_mainSig[2:0] != 3'h0; // @[MulAddRecFN.scala 254:35]
  assign _T_392 = _T_391 | notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 254:39]
  assign notCDom_sig = {notCDom_mainSig[28:3],_T_392}; // @[Cat.scala 30:58]
  assign notCDom_completeCancellation = notCDom_sig[26:25] == 2'h0; // @[MulAddRecFN.scala 257:50]
  assign _T_394 = io_fromPreMul_signProd ^ notCDom_signSigSum; // @[MulAddRecFN.scala 261:36]
  assign notCDom_sign = notCDom_completeCancellation ? roundingMode_min : _T_394; // @[MulAddRecFN.scala 259:12]
  assign notNaN_isInfProd = io_fromPreMul_isInfA | io_fromPreMul_isInfB; // @[MulAddRecFN.scala 266:49]
  assign notNaN_isInfOut = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 267:44]
  assign _T_395 = io_fromPreMul_isZeroA | io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 269:32]
  assign notNaN_addZeros = _T_395 & io_fromPreMul_isZeroC; // @[MulAddRecFN.scala 269:58]
  assign _T_396 = io_fromPreMul_isInfA & io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 274:31]
  assign _T_397 = io_fromPreMul_isSigNaNAny | _T_396; // @[MulAddRecFN.scala 273:35]
  assign _T_398 = io_fromPreMul_isZeroA & io_fromPreMul_isInfB; // @[MulAddRecFN.scala 275:32]
  assign _T_399 = _T_397 | _T_398; // @[MulAddRecFN.scala 274:57]
  assign _T_402 = ~io_fromPreMul_isNaNAOrB & notNaN_isInfProd; // @[MulAddRecFN.scala 276:36]
  assign _T_403 = _T_402 & io_fromPreMul_isInfC; // @[MulAddRecFN.scala 277:61]
  assign _T_404 = _T_403 & io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 278:35]
  assign _T_408 = ~io_fromPreMul_CIsDominant & notCDom_completeCancellation; // @[MulAddRecFN.scala 285:42]
  assign _T_410 = notNaN_isInfProd & io_fromPreMul_signProd; // @[MulAddRecFN.scala 287:27]
  assign _T_411 = io_fromPreMul_isInfC & CDom_sign; // @[MulAddRecFN.scala 288:31]
  assign _T_412 = _T_410 | _T_411; // @[MulAddRecFN.scala 287:54]
  assign _T_414 = notNaN_addZeros & ~roundingMode_min; // @[MulAddRecFN.scala 289:26]
  assign _T_415 = _T_414 & io_fromPreMul_signProd; // @[MulAddRecFN.scala 289:48]
  assign _T_416 = _T_415 & CDom_sign; // @[MulAddRecFN.scala 290:36]
  assign _T_417 = _T_412 | _T_416; // @[MulAddRecFN.scala 288:43]
  assign _T_418 = notNaN_addZeros & roundingMode_min; // @[MulAddRecFN.scala 291:26]
  assign _T_419 = io_fromPreMul_signProd | CDom_sign; // @[MulAddRecFN.scala 292:37]
  assign _T_420 = _T_418 & _T_419; // @[MulAddRecFN.scala 291:46]
  assign _T_421 = _T_417 | _T_420; // @[MulAddRecFN.scala 290:48]
  assign _T_424 = ~notNaN_isInfOut & ~notNaN_addZeros; // @[MulAddRecFN.scala 293:28]
  assign _T_425 = io_fromPreMul_CIsDominant ? CDom_sign : notCDom_sign; // @[MulAddRecFN.scala 294:17]
  assign _T_426 = _T_424 & _T_425; // @[MulAddRecFN.scala 293:49]
  assign io_invalidExc = _T_399 | _T_404; // @[MulAddRecFN.scala 272:19]
  assign io_rawOut_isNaN = io_fromPreMul_isNaNAOrB | io_fromPreMul_isNaNC; // @[MulAddRecFN.scala 280:21]
  assign io_rawOut_isInf = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 281:21]
  assign io_rawOut_isZero = notNaN_addZeros | _T_408; // @[MulAddRecFN.scala 283:22]
  assign io_rawOut_sign = _T_421 | _T_426; // @[MulAddRecFN.scala 286:20]
  assign io_rawOut_sExp = io_fromPreMul_CIsDominant ? $signed(CDom_sExp) : $signed(notCDom_sExp); // @[MulAddRecFN.scala 295:20]
  assign io_rawOut_sig = io_fromPreMul_CIsDominant ? CDom_sig : notCDom_sig; // @[MulAddRecFN.scala 296:19]
  assign MulAddRecFNToRaw_postMul_covSum = 30'h0;
  assign io_covSum = MulAddRecFNToRaw_postMul_covSum;
  assign metaAssert = 1'h0;
endmodule
module RoundAnyRawFNToRecFN_1(
  input         io_in_isZero,
  input         io_in_sign,
  input  [7:0]  io_in_sExp,
  input  [64:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire  _T_11; // @[RoundAnyRawFNToRecFN.scala 96:27]
  wire  _T_13; // @[RoundAnyRawFNToRecFN.scala 96:63]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42]
  wire [8:0] _GEN_0; // @[RoundAnyRawFNToRecFN.scala 102:25]
  wire [9:0] _T_14; // @[RoundAnyRawFNToRecFN.scala 102:25]
  wire [9:0] sAdjustedExp; // @[RoundAnyRawFNToRecFN.scala 104:31]
  wire  _T_18; // @[RoundAnyRawFNToRecFN.scala 115:60]
  wire [26:0] adjustedSig; // @[Cat.scala 30:58]
  wire [26:0] _T_31; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  _T_32; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [26:0] _T_33; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  _T_34; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  common_inexact; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire  _T_36; // @[RoundAnyRawFNToRecFN.scala 167:38]
  wire  _T_37; // @[RoundAnyRawFNToRecFN.scala 167:67]
  wire  _T_38; // @[RoundAnyRawFNToRecFN.scala 169:29]
  wire  _T_39; // @[RoundAnyRawFNToRecFN.scala 168:31]
  wire [26:0] _T_40; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [25:0] _T_42; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _T_43; // @[RoundAnyRawFNToRecFN.scala 173:49]
  wire  _T_45; // @[RoundAnyRawFNToRecFN.scala 173:64]
  wire [25:0] _T_47; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [25:0] _T_49; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [26:0] _T_51; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire  _T_53; // @[RoundAnyRawFNToRecFN.scala 179:42]
  wire [25:0] _T_55; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [25:0] _GEN_1; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] _T_56; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] _T_57; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _T_59; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [9:0] _GEN_2; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [10:0] _T_60; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [8:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [22:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 189:27]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:64]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  wire [8:0] _T_92; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [8:0] expOut; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [22:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [9:0] _T_118; // @[Cat.scala 30:58]
  wire [1:0] _T_120; // @[Cat.scala 30:58]
  wire [29:0] RoundAnyRawFNToRecFN_1_covSum;
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53]
  assign roundingMode_odd = io_roundingMode == 3'h5; // @[RoundAnyRawFNToRecFN.scala 93:53]
  assign _T_11 = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27]
  assign _T_13 = roundingMode_max & ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:63]
  assign roundMagUp = _T_11 | _T_13; // @[RoundAnyRawFNToRecFN.scala 96:42]
  assign _GEN_0 = {{1{io_in_sExp[7]}},io_in_sExp}; // @[RoundAnyRawFNToRecFN.scala 102:25]
  assign _T_14 = $signed(_GEN_0) + 9'shc0; // @[RoundAnyRawFNToRecFN.scala 102:25]
  assign sAdjustedExp = {1'b0,$signed(_T_14[8:0])}; // @[RoundAnyRawFNToRecFN.scala 104:31]
  assign _T_18 = io_in_sig[38:0] != 39'h0; // @[RoundAnyRawFNToRecFN.scala 115:60]
  assign adjustedSig = {io_in_sig[64:39],_T_18}; // @[Cat.scala 30:58]
  assign _T_31 = adjustedSig & 27'h2; // @[RoundAnyRawFNToRecFN.scala 162:40]
  assign _T_32 = _T_31 != 27'h0; // @[RoundAnyRawFNToRecFN.scala 162:56]
  assign _T_33 = adjustedSig & 27'h1; // @[RoundAnyRawFNToRecFN.scala 163:42]
  assign _T_34 = _T_33 != 27'h0; // @[RoundAnyRawFNToRecFN.scala 163:62]
  assign common_inexact = _T_32 | _T_34; // @[RoundAnyRawFNToRecFN.scala 164:36]
  assign _T_36 = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38]
  assign _T_37 = _T_36 & _T_32; // @[RoundAnyRawFNToRecFN.scala 167:67]
  assign _T_38 = roundMagUp & common_inexact; // @[RoundAnyRawFNToRecFN.scala 169:29]
  assign _T_39 = _T_37 | _T_38; // @[RoundAnyRawFNToRecFN.scala 168:31]
  assign _T_40 = adjustedSig | 27'h3; // @[RoundAnyRawFNToRecFN.scala 172:32]
  assign _T_42 = _T_40[26:2] + 25'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  assign _T_43 = roundingMode_near_even & _T_32; // @[RoundAnyRawFNToRecFN.scala 173:49]
  assign _T_45 = _T_43 & ~_T_34; // @[RoundAnyRawFNToRecFN.scala 173:64]
  assign _T_47 = _T_45 ? 26'h1 : 26'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  assign _T_49 = _T_42 & ~_T_47; // @[RoundAnyRawFNToRecFN.scala 172:61]
  assign _T_51 = adjustedSig & 27'h7fffffc; // @[RoundAnyRawFNToRecFN.scala 178:30]
  assign _T_53 = roundingMode_odd & common_inexact; // @[RoundAnyRawFNToRecFN.scala 179:42]
  assign _T_55 = _T_53 ? 26'h1 : 26'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  assign _GEN_1 = {{1'd0}, _T_51[26:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_56 = _GEN_1 | _T_55; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_57 = _T_39 ? _T_49 : _T_56; // @[RoundAnyRawFNToRecFN.scala 171:16]
  assign _T_59 = {1'b0,$signed(_T_57[25:24])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  assign _GEN_2 = {{7{_T_59[2]}},_T_59}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign _T_60 = $signed(sAdjustedExp) + $signed(_GEN_2); // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign common_expOut = _T_60[8:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  assign common_fractOut = _T_57[22:0]; // @[RoundAnyRawFNToRecFN.scala 189:27]
  assign commonCase = ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:64]
  assign inexact = commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  assign _T_92 = io_in_isZero ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign expOut = common_expOut & ~_T_92; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign fractOut = io_in_isZero ? 23'h0 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign _T_118 = {io_in_sign,expOut}; // @[Cat.scala 30:58]
  assign _T_120 = {1'h0,inexact}; // @[Cat.scala 30:58]
  assign io_out = {_T_118,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
  assign io_exceptionFlags = {3'h0,_T_120}; // @[RoundAnyRawFNToRecFN.scala 285:23]
  assign RoundAnyRawFNToRecFN_1_covSum = 30'h0;
  assign io_covSum = RoundAnyRawFNToRecFN_1_covSum;
  assign metaAssert = 1'h0;
endmodule
module RoundAnyRawFNToRecFN_2(
  input         io_in_isZero,
  input         io_in_sign,
  input  [7:0]  io_in_sExp,
  input  [64:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire  _T_11; // @[RoundAnyRawFNToRecFN.scala 96:27]
  wire  _T_13; // @[RoundAnyRawFNToRecFN.scala 96:63]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42]
  wire [11:0] _GEN_0; // @[RoundAnyRawFNToRecFN.scala 102:25]
  wire [12:0] _T_14; // @[RoundAnyRawFNToRecFN.scala 102:25]
  wire [12:0] sAdjustedExp; // @[RoundAnyRawFNToRecFN.scala 104:31]
  wire  _T_18; // @[RoundAnyRawFNToRecFN.scala 115:60]
  wire [55:0] adjustedSig; // @[Cat.scala 30:58]
  wire [55:0] _T_31; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  _T_32; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [55:0] _T_33; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  _T_34; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  common_inexact; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire  _T_36; // @[RoundAnyRawFNToRecFN.scala 167:38]
  wire  _T_37; // @[RoundAnyRawFNToRecFN.scala 167:67]
  wire  _T_38; // @[RoundAnyRawFNToRecFN.scala 169:29]
  wire  _T_39; // @[RoundAnyRawFNToRecFN.scala 168:31]
  wire [55:0] _T_40; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [54:0] _T_42; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _T_43; // @[RoundAnyRawFNToRecFN.scala 173:49]
  wire  _T_45; // @[RoundAnyRawFNToRecFN.scala 173:64]
  wire [54:0] _T_47; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [54:0] _T_49; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [55:0] _T_51; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire  _T_53; // @[RoundAnyRawFNToRecFN.scala 179:42]
  wire [54:0] _T_55; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [54:0] _GEN_1; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [54:0] _T_56; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [54:0] _T_57; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _T_59; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [12:0] _GEN_2; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [13:0] _T_60; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [11:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [51:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 189:27]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:64]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  wire [11:0] _T_92; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [11:0] expOut; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [51:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [12:0] _T_118; // @[Cat.scala 30:58]
  wire [1:0] _T_120; // @[Cat.scala 30:58]
  wire [29:0] RoundAnyRawFNToRecFN_2_covSum;
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53]
  assign roundingMode_odd = io_roundingMode == 3'h5; // @[RoundAnyRawFNToRecFN.scala 93:53]
  assign _T_11 = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27]
  assign _T_13 = roundingMode_max & ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:63]
  assign roundMagUp = _T_11 | _T_13; // @[RoundAnyRawFNToRecFN.scala 96:42]
  assign _GEN_0 = {{4{io_in_sExp[7]}},io_in_sExp}; // @[RoundAnyRawFNToRecFN.scala 102:25]
  assign _T_14 = $signed(_GEN_0) + 12'sh7c0; // @[RoundAnyRawFNToRecFN.scala 102:25]
  assign sAdjustedExp = {1'b0,$signed(_T_14[11:0])}; // @[RoundAnyRawFNToRecFN.scala 104:31]
  assign _T_18 = io_in_sig[9:0] != 10'h0; // @[RoundAnyRawFNToRecFN.scala 115:60]
  assign adjustedSig = {io_in_sig[64:10],_T_18}; // @[Cat.scala 30:58]
  assign _T_31 = adjustedSig & 56'h2; // @[RoundAnyRawFNToRecFN.scala 162:40]
  assign _T_32 = _T_31 != 56'h0; // @[RoundAnyRawFNToRecFN.scala 162:56]
  assign _T_33 = adjustedSig & 56'h1; // @[RoundAnyRawFNToRecFN.scala 163:42]
  assign _T_34 = _T_33 != 56'h0; // @[RoundAnyRawFNToRecFN.scala 163:62]
  assign common_inexact = _T_32 | _T_34; // @[RoundAnyRawFNToRecFN.scala 164:36]
  assign _T_36 = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38]
  assign _T_37 = _T_36 & _T_32; // @[RoundAnyRawFNToRecFN.scala 167:67]
  assign _T_38 = roundMagUp & common_inexact; // @[RoundAnyRawFNToRecFN.scala 169:29]
  assign _T_39 = _T_37 | _T_38; // @[RoundAnyRawFNToRecFN.scala 168:31]
  assign _T_40 = adjustedSig | 56'h3; // @[RoundAnyRawFNToRecFN.scala 172:32]
  assign _T_42 = _T_40[55:2] + 54'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  assign _T_43 = roundingMode_near_even & _T_32; // @[RoundAnyRawFNToRecFN.scala 173:49]
  assign _T_45 = _T_43 & ~_T_34; // @[RoundAnyRawFNToRecFN.scala 173:64]
  assign _T_47 = _T_45 ? 55'h1 : 55'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  assign _T_49 = _T_42 & ~_T_47; // @[RoundAnyRawFNToRecFN.scala 172:61]
  assign _T_51 = adjustedSig & 56'hfffffffffffffc; // @[RoundAnyRawFNToRecFN.scala 178:30]
  assign _T_53 = roundingMode_odd & common_inexact; // @[RoundAnyRawFNToRecFN.scala 179:42]
  assign _T_55 = _T_53 ? 55'h1 : 55'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  assign _GEN_1 = {{1'd0}, _T_51[55:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_56 = _GEN_1 | _T_55; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_57 = _T_39 ? _T_49 : _T_56; // @[RoundAnyRawFNToRecFN.scala 171:16]
  assign _T_59 = {1'b0,$signed(_T_57[54:53])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  assign _GEN_2 = {{10{_T_59[2]}},_T_59}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign _T_60 = $signed(sAdjustedExp) + $signed(_GEN_2); // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign common_expOut = _T_60[11:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  assign common_fractOut = _T_57[51:0]; // @[RoundAnyRawFNToRecFN.scala 189:27]
  assign commonCase = ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:64]
  assign inexact = commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  assign _T_92 = io_in_isZero ? 12'he00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign expOut = common_expOut & ~_T_92; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign fractOut = io_in_isZero ? 52'h0 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign _T_118 = {io_in_sign,expOut}; // @[Cat.scala 30:58]
  assign _T_120 = {1'h0,inexact}; // @[Cat.scala 30:58]
  assign io_out = {_T_118,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
  assign io_exceptionFlags = {3'h0,_T_120}; // @[RoundAnyRawFNToRecFN.scala 285:23]
  assign RoundAnyRawFNToRecFN_2_covSum = 30'h0;
  assign io_covSum = RoundAnyRawFNToRecFN_2_covSum;
  assign metaAssert = 1'h0;
endmodule
module RoundAnyRawFNToRecFN_3(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [12:0] io_in_sExp,
  input  [53:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire  _T_11; // @[RoundAnyRawFNToRecFN.scala 96:27]
  wire  _T_13; // @[RoundAnyRawFNToRecFN.scala 96:63]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42]
  wire [13:0] sAdjustedExp; // @[RoundAnyRawFNToRecFN.scala 108:24]
  wire  _T_16; // @[RoundAnyRawFNToRecFN.scala 115:60]
  wire [26:0] adjustedSig; // @[Cat.scala 30:58]
  wire  _T_25; // @[primitives.scala 57:25]
  wire  _T_27; // @[primitives.scala 57:25]
  wire  _T_29; // @[primitives.scala 57:25]
  wire [5:0] _T_30; // @[primitives.scala 58:26]
  wire [64:0] _T_31; // @[primitives.scala 77:58]
  wire [15:0] _T_37; // @[Bitwise.scala 103:31]
  wire [15:0] _T_39; // @[Bitwise.scala 103:65]
  wire [15:0] _T_41; // @[Bitwise.scala 103:75]
  wire [15:0] _T_42; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_0; // @[Bitwise.scala 103:31]
  wire [15:0] _T_47; // @[Bitwise.scala 103:31]
  wire [15:0] _T_49; // @[Bitwise.scala 103:65]
  wire [15:0] _T_51; // @[Bitwise.scala 103:75]
  wire [15:0] _T_52; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_1; // @[Bitwise.scala 103:31]
  wire [15:0] _T_57; // @[Bitwise.scala 103:31]
  wire [15:0] _T_59; // @[Bitwise.scala 103:65]
  wire [15:0] _T_61; // @[Bitwise.scala 103:75]
  wire [15:0] _T_62; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_2; // @[Bitwise.scala 103:31]
  wire [15:0] _T_67; // @[Bitwise.scala 103:31]
  wire [15:0] _T_69; // @[Bitwise.scala 103:65]
  wire [15:0] _T_71; // @[Bitwise.scala 103:75]
  wire [15:0] _T_72; // @[Bitwise.scala 103:39]
  wire [21:0] _T_89; // @[Cat.scala 30:58]
  wire [21:0] _T_91; // @[primitives.scala 74:21]
  wire [24:0] _T_93; // @[Cat.scala 30:58]
  wire [2:0] _T_103; // @[Cat.scala 30:58]
  wire [2:0] _T_104; // @[primitives.scala 61:24]
  wire [24:0] _T_105; // @[primitives.scala 66:24]
  wire [24:0] _T_106; // @[primitives.scala 61:24]
  wire [26:0] _T_108; // @[Cat.scala 30:58]
  wire [26:0] _T_110; // @[Cat.scala 30:58]
  wire [26:0] _T_112; // @[RoundAnyRawFNToRecFN.scala 161:46]
  wire [26:0] _T_113; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  _T_114; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [26:0] _T_115; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  _T_116; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  _T_117; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire  _T_118; // @[RoundAnyRawFNToRecFN.scala 167:38]
  wire  _T_119; // @[RoundAnyRawFNToRecFN.scala 167:67]
  wire  _T_120; // @[RoundAnyRawFNToRecFN.scala 169:29]
  wire  _T_121; // @[RoundAnyRawFNToRecFN.scala 168:31]
  wire [26:0] _T_122; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [25:0] _T_124; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _T_125; // @[RoundAnyRawFNToRecFN.scala 173:49]
  wire  _T_127; // @[RoundAnyRawFNToRecFN.scala 173:64]
  wire [25:0] _T_129; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [25:0] _T_131; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [26:0] _T_133; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire  _T_135; // @[RoundAnyRawFNToRecFN.scala 179:42]
  wire [25:0] _T_137; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [25:0] _GEN_3; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] _T_138; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] _T_139; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _T_141; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [13:0] _GEN_4; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [14:0] _T_142; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [8:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [22:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 189:27]
  wire [7:0] _T_147; // @[RoundAnyRawFNToRecFN.scala 194:30]
  wire  common_overflow; // @[RoundAnyRawFNToRecFN.scala 194:50]
  wire  common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 198:31]
  wire  _T_156; // @[RoundAnyRawFNToRecFN.scala 203:70]
  wire  _T_159; // @[RoundAnyRawFNToRecFN.scala 205:67]
  wire  _T_160; // @[RoundAnyRawFNToRecFN.scala 207:29]
  wire  _T_161; // @[RoundAnyRawFNToRecFN.scala 206:46]
  wire [5:0] _T_165; // @[RoundAnyRawFNToRecFN.scala 218:48]
  wire  _T_166; // @[RoundAnyRawFNToRecFN.scala 218:62]
  wire  _T_167; // @[RoundAnyRawFNToRecFN.scala 218:32]
  wire  _T_171; // @[RoundAnyRawFNToRecFN.scala 218:74]
  wire  _T_178; // @[RoundAnyRawFNToRecFN.scala 224:38]
  wire  _T_179; // @[RoundAnyRawFNToRecFN.scala 225:45]
  wire  _T_180; // @[RoundAnyRawFNToRecFN.scala 225:60]
  wire  _T_182; // @[RoundAnyRawFNToRecFN.scala 219:76]
  wire  common_underflow; // @[RoundAnyRawFNToRecFN.scala 215:40]
  wire  common_inexact; // @[RoundAnyRawFNToRecFN.scala 228:49]
  wire  isNaNOut; // @[RoundAnyRawFNToRecFN.scala 233:34]
  wire  _T_187; // @[RoundAnyRawFNToRecFN.scala 235:33]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:61]
  wire  overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  wire  underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  wire  _T_189; // @[RoundAnyRawFNToRecFN.scala 238:43]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:28]
  wire  overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  wire  _T_191; // @[RoundAnyRawFNToRecFN.scala 243:20]
  wire  _T_192; // @[RoundAnyRawFNToRecFN.scala 243:60]
  wire  pegMinNonzeroMagOut; // @[RoundAnyRawFNToRecFN.scala 243:45]
  wire  pegMaxFiniteMagOut; // @[RoundAnyRawFNToRecFN.scala 244:39]
  wire  _T_194; // @[RoundAnyRawFNToRecFN.scala 246:45]
  wire  notNaN_isInfOut; // @[RoundAnyRawFNToRecFN.scala 246:32]
  wire  signOut; // @[RoundAnyRawFNToRecFN.scala 248:22]
  wire  _T_195; // @[RoundAnyRawFNToRecFN.scala 251:32]
  wire [8:0] _T_196; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [8:0] _T_198; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [8:0] _T_200; // @[RoundAnyRawFNToRecFN.scala 255:18]
  wire [8:0] _T_202; // @[RoundAnyRawFNToRecFN.scala 254:17]
  wire [8:0] _T_203; // @[RoundAnyRawFNToRecFN.scala 259:18]
  wire [8:0] _T_205; // @[RoundAnyRawFNToRecFN.scala 258:17]
  wire [8:0] _T_206; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [8:0] _T_208; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [8:0] _T_209; // @[RoundAnyRawFNToRecFN.scala 267:16]
  wire [8:0] _T_210; // @[RoundAnyRawFNToRecFN.scala 266:18]
  wire [8:0] _T_211; // @[RoundAnyRawFNToRecFN.scala 271:16]
  wire [8:0] _T_212; // @[RoundAnyRawFNToRecFN.scala 270:15]
  wire [8:0] _T_213; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [8:0] _T_214; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [8:0] _T_215; // @[RoundAnyRawFNToRecFN.scala 276:16]
  wire [8:0] expOut; // @[RoundAnyRawFNToRecFN.scala 275:77]
  wire  _T_216; // @[RoundAnyRawFNToRecFN.scala 278:22]
  wire  _T_217; // @[RoundAnyRawFNToRecFN.scala 278:38]
  wire [22:0] _T_218; // @[RoundAnyRawFNToRecFN.scala 279:16]
  wire [22:0] _T_219; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [22:0] _T_221; // @[Bitwise.scala 72:12]
  wire [22:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 281:11]
  wire [9:0] _T_222; // @[Cat.scala 30:58]
  wire [1:0] _T_224; // @[Cat.scala 30:58]
  wire [2:0] _T_226; // @[Cat.scala 30:58]
  wire [29:0] RoundAnyRawFNToRecFN_3_covSum;
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53]
  assign roundingMode_odd = io_roundingMode == 3'h5; // @[RoundAnyRawFNToRecFN.scala 93:53]
  assign _T_11 = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27]
  assign _T_13 = roundingMode_max & ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:63]
  assign roundMagUp = _T_11 | _T_13; // @[RoundAnyRawFNToRecFN.scala 96:42]
  assign sAdjustedExp = $signed(io_in_sExp) + -13'sh700; // @[RoundAnyRawFNToRecFN.scala 108:24]
  assign _T_16 = io_in_sig[27:0] != 28'h0; // @[RoundAnyRawFNToRecFN.scala 115:60]
  assign adjustedSig = {io_in_sig[53:28],_T_16}; // @[Cat.scala 30:58]
  assign _T_25 = ~sAdjustedExp[8]; // @[primitives.scala 57:25]
  assign _T_27 = ~sAdjustedExp[7]; // @[primitives.scala 57:25]
  assign _T_29 = ~sAdjustedExp[6]; // @[primitives.scala 57:25]
  assign _T_30 = ~sAdjustedExp[5:0]; // @[primitives.scala 58:26]
  assign _T_31 = -65'sh10000000000000000 >>> _T_30; // @[primitives.scala 77:58]
  assign _T_37 = {{8'd0}, _T_31[57:50]}; // @[Bitwise.scala 103:31]
  assign _T_39 = {_T_31[49:42], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_41 = _T_39 & 16'hff00; // @[Bitwise.scala 103:75]
  assign _T_42 = _T_37 | _T_41; // @[Bitwise.scala 103:39]
  assign _GEN_0 = {{4'd0}, _T_42[15:4]}; // @[Bitwise.scala 103:31]
  assign _T_47 = _GEN_0 & 16'hf0f; // @[Bitwise.scala 103:31]
  assign _T_49 = {_T_42[11:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_51 = _T_49 & 16'hf0f0; // @[Bitwise.scala 103:75]
  assign _T_52 = _T_47 | _T_51; // @[Bitwise.scala 103:39]
  assign _GEN_1 = {{2'd0}, _T_52[15:2]}; // @[Bitwise.scala 103:31]
  assign _T_57 = _GEN_1 & 16'h3333; // @[Bitwise.scala 103:31]
  assign _T_59 = {_T_52[13:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_61 = _T_59 & 16'hcccc; // @[Bitwise.scala 103:75]
  assign _T_62 = _T_57 | _T_61; // @[Bitwise.scala 103:39]
  assign _GEN_2 = {{1'd0}, _T_62[15:1]}; // @[Bitwise.scala 103:31]
  assign _T_67 = _GEN_2 & 16'h5555; // @[Bitwise.scala 103:31]
  assign _T_69 = {_T_62[14:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_71 = _T_69 & 16'haaaa; // @[Bitwise.scala 103:75]
  assign _T_72 = _T_67 | _T_71; // @[Bitwise.scala 103:39]
  assign _T_89 = {_T_72,_T_31[58],_T_31[59],_T_31[60],_T_31[61],_T_31[62],_T_31[63]}; // @[Cat.scala 30:58]
  assign _T_91 = _T_29 ? 22'h0 : ~_T_89; // @[primitives.scala 74:21]
  assign _T_93 = {~_T_91,3'h7}; // @[Cat.scala 30:58]
  assign _T_103 = {_T_31[0],_T_31[1],_T_31[2]}; // @[Cat.scala 30:58]
  assign _T_104 = _T_29 ? _T_103 : 3'h0; // @[primitives.scala 61:24]
  assign _T_105 = _T_27 ? _T_93 : {{22'd0}, _T_104}; // @[primitives.scala 66:24]
  assign _T_106 = _T_25 ? _T_105 : 25'h0; // @[primitives.scala 61:24]
  assign _T_108 = {_T_106,2'h3}; // @[Cat.scala 30:58]
  assign _T_110 = {1'h0,_T_108[26:1]}; // @[Cat.scala 30:58]
  assign _T_112 = ~_T_110 & _T_108; // @[RoundAnyRawFNToRecFN.scala 161:46]
  assign _T_113 = adjustedSig & _T_112; // @[RoundAnyRawFNToRecFN.scala 162:40]
  assign _T_114 = _T_113 != 27'h0; // @[RoundAnyRawFNToRecFN.scala 162:56]
  assign _T_115 = adjustedSig & _T_110; // @[RoundAnyRawFNToRecFN.scala 163:42]
  assign _T_116 = _T_115 != 27'h0; // @[RoundAnyRawFNToRecFN.scala 163:62]
  assign _T_117 = _T_114 | _T_116; // @[RoundAnyRawFNToRecFN.scala 164:36]
  assign _T_118 = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38]
  assign _T_119 = _T_118 & _T_114; // @[RoundAnyRawFNToRecFN.scala 167:67]
  assign _T_120 = roundMagUp & _T_117; // @[RoundAnyRawFNToRecFN.scala 169:29]
  assign _T_121 = _T_119 | _T_120; // @[RoundAnyRawFNToRecFN.scala 168:31]
  assign _T_122 = adjustedSig | _T_108; // @[RoundAnyRawFNToRecFN.scala 172:32]
  assign _T_124 = _T_122[26:2] + 25'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  assign _T_125 = roundingMode_near_even & _T_114; // @[RoundAnyRawFNToRecFN.scala 173:49]
  assign _T_127 = _T_125 & ~_T_116; // @[RoundAnyRawFNToRecFN.scala 173:64]
  assign _T_129 = _T_127 ? _T_108[26:1] : 26'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  assign _T_131 = _T_124 & ~_T_129; // @[RoundAnyRawFNToRecFN.scala 172:61]
  assign _T_133 = adjustedSig & ~_T_108; // @[RoundAnyRawFNToRecFN.scala 178:30]
  assign _T_135 = roundingMode_odd & _T_117; // @[RoundAnyRawFNToRecFN.scala 179:42]
  assign _T_137 = _T_135 ? _T_112[26:1] : 26'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  assign _GEN_3 = {{1'd0}, _T_133[26:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_138 = _GEN_3 | _T_137; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_139 = _T_121 ? _T_131 : _T_138; // @[RoundAnyRawFNToRecFN.scala 171:16]
  assign _T_141 = {1'b0,$signed(_T_139[25:24])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  assign _GEN_4 = {{11{_T_141[2]}},_T_141}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign _T_142 = $signed(sAdjustedExp) + $signed(_GEN_4); // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign common_expOut = _T_142[8:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  assign common_fractOut = _T_139[22:0]; // @[RoundAnyRawFNToRecFN.scala 189:27]
  assign _T_147 = _T_142[14:7]; // @[RoundAnyRawFNToRecFN.scala 194:30]
  assign common_overflow = $signed(_T_147) >= 8'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50]
  assign common_totalUnderflow = $signed(_T_142) < 15'sh6b; // @[RoundAnyRawFNToRecFN.scala 198:31]
  assign _T_156 = adjustedSig[1:0] != 2'h0; // @[RoundAnyRawFNToRecFN.scala 203:70]
  assign _T_159 = _T_118 & adjustedSig[1]; // @[RoundAnyRawFNToRecFN.scala 205:67]
  assign _T_160 = roundMagUp & _T_156; // @[RoundAnyRawFNToRecFN.scala 207:29]
  assign _T_161 = _T_159 | _T_160; // @[RoundAnyRawFNToRecFN.scala 206:46]
  assign _T_165 = sAdjustedExp[13:8]; // @[RoundAnyRawFNToRecFN.scala 218:48]
  assign _T_166 = $signed(_T_165) <= 6'sh0; // @[RoundAnyRawFNToRecFN.scala 218:62]
  assign _T_167 = _T_117 & _T_166; // @[RoundAnyRawFNToRecFN.scala 218:32]
  assign _T_171 = _T_167 & _T_108[2]; // @[RoundAnyRawFNToRecFN.scala 218:74]
  assign _T_178 = ~_T_108[3] & _T_139[24]; // @[RoundAnyRawFNToRecFN.scala 224:38]
  assign _T_179 = _T_178 & _T_114; // @[RoundAnyRawFNToRecFN.scala 225:45]
  assign _T_180 = _T_179 & _T_161; // @[RoundAnyRawFNToRecFN.scala 225:60]
  assign _T_182 = _T_171 & ~_T_180; // @[RoundAnyRawFNToRecFN.scala 219:76]
  assign common_underflow = common_totalUnderflow | _T_182; // @[RoundAnyRawFNToRecFN.scala 215:40]
  assign common_inexact = common_totalUnderflow | _T_117; // @[RoundAnyRawFNToRecFN.scala 228:49]
  assign isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34]
  assign _T_187 = ~isNaNOut & ~io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 235:33]
  assign commonCase = _T_187 & ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:61]
  assign overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  assign underflow = commonCase & common_underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  assign _T_189 = commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  assign inexact = overflow | _T_189; // @[RoundAnyRawFNToRecFN.scala 238:28]
  assign overflow_roundMagUp = _T_118 | roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  assign _T_191 = commonCase & common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 243:20]
  assign _T_192 = roundMagUp | roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 243:60]
  assign pegMinNonzeroMagOut = _T_191 & _T_192; // @[RoundAnyRawFNToRecFN.scala 243:45]
  assign pegMaxFiniteMagOut = overflow & ~overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 244:39]
  assign _T_194 = overflow & overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 246:45]
  assign notNaN_isInfOut = io_in_isInf | _T_194; // @[RoundAnyRawFNToRecFN.scala 246:32]
  assign signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22]
  assign _T_195 = io_in_isZero | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 251:32]
  assign _T_196 = _T_195 ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign _T_198 = common_expOut & ~_T_196; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign _T_200 = pegMinNonzeroMagOut ? 9'h194 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 255:18]
  assign _T_202 = _T_198 & ~_T_200; // @[RoundAnyRawFNToRecFN.scala 254:17]
  assign _T_203 = pegMaxFiniteMagOut ? 9'h80 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 259:18]
  assign _T_205 = _T_202 & ~_T_203; // @[RoundAnyRawFNToRecFN.scala 258:17]
  assign _T_206 = notNaN_isInfOut ? 9'h40 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  assign _T_208 = _T_205 & ~_T_206; // @[RoundAnyRawFNToRecFN.scala 262:17]
  assign _T_209 = pegMinNonzeroMagOut ? 9'h6b : 9'h0; // @[RoundAnyRawFNToRecFN.scala 267:16]
  assign _T_210 = _T_208 | _T_209; // @[RoundAnyRawFNToRecFN.scala 266:18]
  assign _T_211 = pegMaxFiniteMagOut ? 9'h17f : 9'h0; // @[RoundAnyRawFNToRecFN.scala 271:16]
  assign _T_212 = _T_210 | _T_211; // @[RoundAnyRawFNToRecFN.scala 270:15]
  assign _T_213 = notNaN_isInfOut ? 9'h180 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  assign _T_214 = _T_212 | _T_213; // @[RoundAnyRawFNToRecFN.scala 274:15]
  assign _T_215 = isNaNOut ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 276:16]
  assign expOut = _T_214 | _T_215; // @[RoundAnyRawFNToRecFN.scala 275:77]
  assign _T_216 = isNaNOut | io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 278:22]
  assign _T_217 = _T_216 | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 278:38]
  assign _T_218 = isNaNOut ? 23'h400000 : 23'h0; // @[RoundAnyRawFNToRecFN.scala 279:16]
  assign _T_219 = _T_217 ? _T_218 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign _T_221 = pegMaxFiniteMagOut ? 23'h7fffff : 23'h0; // @[Bitwise.scala 72:12]
  assign fractOut = _T_219 | _T_221; // @[RoundAnyRawFNToRecFN.scala 281:11]
  assign _T_222 = {signOut,expOut}; // @[Cat.scala 30:58]
  assign _T_224 = {underflow,inexact}; // @[Cat.scala 30:58]
  assign _T_226 = {io_invalidExc,1'h0,overflow}; // @[Cat.scala 30:58]
  assign io_out = {_T_222,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
  assign io_exceptionFlags = {_T_226,_T_224}; // @[RoundAnyRawFNToRecFN.scala 285:23]
  assign RoundAnyRawFNToRecFN_3_covSum = 30'h0;
  assign io_covSum = RoundAnyRawFNToRecFN_3_covSum;
  assign metaAssert = 1'h0;
endmodule
module MulAddRecFNToRaw_preMul_1(
  input  [1:0]   io_op,
  input  [64:0]  io_a,
  input  [64:0]  io_b,
  input  [64:0]  io_c,
  output [52:0]  io_mulAddA,
  output [52:0]  io_mulAddB,
  output [105:0] io_mulAddC,
  output         io_toPostMul_isSigNaNAny,
  output         io_toPostMul_isNaNAOrB,
  output         io_toPostMul_isInfA,
  output         io_toPostMul_isZeroA,
  output         io_toPostMul_isInfB,
  output         io_toPostMul_isZeroB,
  output         io_toPostMul_signProd,
  output         io_toPostMul_isNaNC,
  output         io_toPostMul_isInfC,
  output         io_toPostMul_isZeroC,
  output [12:0]  io_toPostMul_sExpSum,
  output         io_toPostMul_doSubMags,
  output         io_toPostMul_CIsDominant,
  output [5:0]   io_toPostMul_CDom_CAlignDist,
  output [54:0]  io_toPostMul_highAlignedSigC,
  output         io_toPostMul_bit0AlignedSigC,
  output [29:0]  io_covSum,
  output         metaAssert
);
  wire  rawA_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_16; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawA_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawA_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] rawA_sig; // @[Cat.scala 30:58]
  wire  rawB_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_33; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawB_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawB_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] rawB_sig; // @[Cat.scala 30:58]
  wire  rawC_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_50; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawC_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawC_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawC_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] rawC_sig; // @[Cat.scala 30:58]
  wire  _T_63; // @[MulAddRecFN.scala 98:30]
  wire  signProd; // @[MulAddRecFN.scala 98:42]
  wire [13:0] _T_65; // @[MulAddRecFN.scala 101:19]
  wire [13:0] sExpAlignedProd; // @[MulAddRecFN.scala 101:32]
  wire  _T_68; // @[MulAddRecFN.scala 103:30]
  wire  doSubMags; // @[MulAddRecFN.scala 103:42]
  wire [13:0] _GEN_0; // @[MulAddRecFN.scala 107:42]
  wire [13:0] sNatCAlignDist; // @[MulAddRecFN.scala 107:42]
  wire [12:0] posNatCAlignDist; // @[MulAddRecFN.scala 108:42]
  wire  _T_72; // @[MulAddRecFN.scala 109:35]
  wire  _T_73; // @[MulAddRecFN.scala 109:69]
  wire  isMinCAlign; // @[MulAddRecFN.scala 109:50]
  wire  _T_75; // @[MulAddRecFN.scala 111:60]
  wire  _T_76; // @[MulAddRecFN.scala 111:39]
  wire  CIsDominant; // @[MulAddRecFN.scala 111:23]
  wire  _T_77; // @[MulAddRecFN.scala 115:34]
  wire [7:0] _T_79; // @[MulAddRecFN.scala 115:16]
  wire [7:0] CAlignDist; // @[MulAddRecFN.scala 113:12]
  wire [53:0] _T_81; // @[MulAddRecFN.scala 121:16]
  wire [110:0] _T_83; // @[Bitwise.scala 72:12]
  wire [164:0] _T_85; // @[MulAddRecFN.scala 123:11]
  wire [164:0] mainAlignedSigC; // @[MulAddRecFN.scala 123:17]
  wire  _T_108; // @[primitives.scala 121:54]
  wire  _T_110; // @[primitives.scala 121:54]
  wire  _T_112; // @[primitives.scala 121:54]
  wire  _T_114; // @[primitives.scala 121:54]
  wire  _T_116; // @[primitives.scala 121:54]
  wire  _T_118; // @[primitives.scala 121:54]
  wire  _T_120; // @[primitives.scala 121:54]
  wire  _T_122; // @[primitives.scala 121:54]
  wire  _T_124; // @[primitives.scala 121:54]
  wire  _T_126; // @[primitives.scala 121:54]
  wire  _T_128; // @[primitives.scala 121:54]
  wire  _T_130; // @[primitives.scala 121:54]
  wire  _T_132; // @[primitives.scala 121:54]
  wire  _T_134; // @[primitives.scala 124:57]
  wire [6:0] _T_140; // @[primitives.scala 125:20]
  wire [13:0] _T_147; // @[primitives.scala 125:20]
  wire [64:0] _T_149; // @[primitives.scala 77:58]
  wire [7:0] _T_155; // @[Bitwise.scala 103:31]
  wire [7:0] _T_157; // @[Bitwise.scala 103:65]
  wire [7:0] _T_159; // @[Bitwise.scala 103:75]
  wire [7:0] _T_160; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_1; // @[Bitwise.scala 103:31]
  wire [7:0] _T_165; // @[Bitwise.scala 103:31]
  wire [7:0] _T_167; // @[Bitwise.scala 103:65]
  wire [7:0] _T_169; // @[Bitwise.scala 103:75]
  wire [7:0] _T_170; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_2; // @[Bitwise.scala 103:31]
  wire [7:0] _T_175; // @[Bitwise.scala 103:31]
  wire [7:0] _T_177; // @[Bitwise.scala 103:65]
  wire [7:0] _T_179; // @[Bitwise.scala 103:75]
  wire [7:0] _T_180; // @[Bitwise.scala 103:39]
  wire [12:0] _T_194; // @[Cat.scala 30:58]
  wire [13:0] _GEN_3; // @[MulAddRecFN.scala 125:68]
  wire [13:0] _T_195; // @[MulAddRecFN.scala 125:68]
  wire  reduced4CExtra; // @[MulAddRecFN.scala 133:11]
  wire  _T_199; // @[MulAddRecFN.scala 137:39]
  wire  _T_201; // @[MulAddRecFN.scala 137:44]
  wire  _T_203; // @[MulAddRecFN.scala 138:39]
  wire  _T_204; // @[MulAddRecFN.scala 138:44]
  wire  _T_205; // @[MulAddRecFN.scala 136:16]
  wire [161:0] _T_206; // @[Cat.scala 30:58]
  wire [162:0] alignedSigC; // @[Cat.scala 30:58]
  wire  _T_210; // @[common.scala 81:46]
  wire  _T_213; // @[common.scala 81:46]
  wire  _T_214; // @[MulAddRecFN.scala 149:32]
  wire  _T_217; // @[common.scala 81:46]
  wire [13:0] _T_222; // @[MulAddRecFN.scala 161:53]
  wire [13:0] _T_223; // @[MulAddRecFN.scala 161:12]
  wire [29:0] MulAddRecFNToRaw_preMul_1_covSum;
  assign rawA_isZero = io_a[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_16 = io_a[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawA_isNaN = _T_16 & io_a[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawA_sign = io_a[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawA_sExp = {1'b0,$signed(io_a[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawA_sig = {1'h0,~rawA_isZero,io_a[51:0]}; // @[Cat.scala 30:58]
  assign rawB_isZero = io_b[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_33 = io_b[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawB_isNaN = _T_33 & io_b[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawB_sign = io_b[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawB_sExp = {1'b0,$signed(io_b[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawB_sig = {1'h0,~rawB_isZero,io_b[51:0]}; // @[Cat.scala 30:58]
  assign rawC_isZero = io_c[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_50 = io_c[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawC_isNaN = _T_50 & io_c[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawC_sign = io_c[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawC_sExp = {1'b0,$signed(io_c[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawC_sig = {1'h0,~rawC_isZero,io_c[51:0]}; // @[Cat.scala 30:58]
  assign _T_63 = rawA_sign ^ rawB_sign; // @[MulAddRecFN.scala 98:30]
  assign signProd = _T_63 ^ io_op[1]; // @[MulAddRecFN.scala 98:42]
  assign _T_65 = $signed(rawA_sExp) + $signed(rawB_sExp); // @[MulAddRecFN.scala 101:19]
  assign sExpAlignedProd = $signed(_T_65) + -14'sh7c8; // @[MulAddRecFN.scala 101:32]
  assign _T_68 = signProd ^ rawC_sign; // @[MulAddRecFN.scala 103:30]
  assign doSubMags = _T_68 ^ io_op[0]; // @[MulAddRecFN.scala 103:42]
  assign _GEN_0 = {{1{rawC_sExp[12]}},rawC_sExp}; // @[MulAddRecFN.scala 107:42]
  assign sNatCAlignDist = $signed(sExpAlignedProd) - $signed(_GEN_0); // @[MulAddRecFN.scala 107:42]
  assign posNatCAlignDist = sNatCAlignDist[12:0]; // @[MulAddRecFN.scala 108:42]
  assign _T_72 = rawA_isZero | rawB_isZero; // @[MulAddRecFN.scala 109:35]
  assign _T_73 = $signed(sNatCAlignDist) < 14'sh0; // @[MulAddRecFN.scala 109:69]
  assign isMinCAlign = _T_72 | _T_73; // @[MulAddRecFN.scala 109:50]
  assign _T_75 = posNatCAlignDist <= 13'h35; // @[MulAddRecFN.scala 111:60]
  assign _T_76 = isMinCAlign | _T_75; // @[MulAddRecFN.scala 111:39]
  assign CIsDominant = ~rawC_isZero & _T_76; // @[MulAddRecFN.scala 111:23]
  assign _T_77 = posNatCAlignDist < 13'ha1; // @[MulAddRecFN.scala 115:34]
  assign _T_79 = _T_77 ? posNatCAlignDist[7:0] : 8'ha1; // @[MulAddRecFN.scala 115:16]
  assign CAlignDist = isMinCAlign ? 8'h0 : _T_79; // @[MulAddRecFN.scala 113:12]
  assign _T_81 = doSubMags ? ~rawC_sig : rawC_sig; // @[MulAddRecFN.scala 121:16]
  assign _T_83 = doSubMags ? 111'h7fffffffffffffffffffffffffff : 111'h0; // @[Bitwise.scala 72:12]
  assign _T_85 = {_T_81,_T_83}; // @[MulAddRecFN.scala 123:11]
  assign mainAlignedSigC = $signed(_T_85) >>> CAlignDist; // @[MulAddRecFN.scala 123:17]
  assign _T_108 = rawC_sig[3:0] != 4'h0; // @[primitives.scala 121:54]
  assign _T_110 = rawC_sig[7:4] != 4'h0; // @[primitives.scala 121:54]
  assign _T_112 = rawC_sig[11:8] != 4'h0; // @[primitives.scala 121:54]
  assign _T_114 = rawC_sig[15:12] != 4'h0; // @[primitives.scala 121:54]
  assign _T_116 = rawC_sig[19:16] != 4'h0; // @[primitives.scala 121:54]
  assign _T_118 = rawC_sig[23:20] != 4'h0; // @[primitives.scala 121:54]
  assign _T_120 = rawC_sig[27:24] != 4'h0; // @[primitives.scala 121:54]
  assign _T_122 = rawC_sig[31:28] != 4'h0; // @[primitives.scala 121:54]
  assign _T_124 = rawC_sig[35:32] != 4'h0; // @[primitives.scala 121:54]
  assign _T_126 = rawC_sig[39:36] != 4'h0; // @[primitives.scala 121:54]
  assign _T_128 = rawC_sig[43:40] != 4'h0; // @[primitives.scala 121:54]
  assign _T_130 = rawC_sig[47:44] != 4'h0; // @[primitives.scala 121:54]
  assign _T_132 = rawC_sig[51:48] != 4'h0; // @[primitives.scala 121:54]
  assign _T_134 = rawC_sig[53:52] != 2'h0; // @[primitives.scala 124:57]
  assign _T_140 = {_T_120,_T_118,_T_116,_T_114,_T_112,_T_110,_T_108}; // @[primitives.scala 125:20]
  assign _T_147 = {_T_134,_T_132,_T_130,_T_128,_T_126,_T_124,_T_122,_T_140}; // @[primitives.scala 125:20]
  assign _T_149 = -65'sh10000000000000000 >>> CAlignDist[7:2]; // @[primitives.scala 77:58]
  assign _T_155 = {{4'd0}, _T_149[31:28]}; // @[Bitwise.scala 103:31]
  assign _T_157 = {_T_149[27:24], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_159 = _T_157 & 8'hf0; // @[Bitwise.scala 103:75]
  assign _T_160 = _T_155 | _T_159; // @[Bitwise.scala 103:39]
  assign _GEN_1 = {{2'd0}, _T_160[7:2]}; // @[Bitwise.scala 103:31]
  assign _T_165 = _GEN_1 & 8'h33; // @[Bitwise.scala 103:31]
  assign _T_167 = {_T_160[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_169 = _T_167 & 8'hcc; // @[Bitwise.scala 103:75]
  assign _T_170 = _T_165 | _T_169; // @[Bitwise.scala 103:39]
  assign _GEN_2 = {{1'd0}, _T_170[7:1]}; // @[Bitwise.scala 103:31]
  assign _T_175 = _GEN_2 & 8'h55; // @[Bitwise.scala 103:31]
  assign _T_177 = {_T_170[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_179 = _T_177 & 8'haa; // @[Bitwise.scala 103:75]
  assign _T_180 = _T_175 | _T_179; // @[Bitwise.scala 103:39]
  assign _T_194 = {_T_180,_T_149[32],_T_149[33],_T_149[34],_T_149[35],_T_149[36]}; // @[Cat.scala 30:58]
  assign _GEN_3 = {{1'd0}, _T_194}; // @[MulAddRecFN.scala 125:68]
  assign _T_195 = _T_147 & _GEN_3; // @[MulAddRecFN.scala 125:68]
  assign reduced4CExtra = _T_195 != 14'h0; // @[MulAddRecFN.scala 133:11]
  assign _T_199 = ~mainAlignedSigC[2:0] == 3'h0; // @[MulAddRecFN.scala 137:39]
  assign _T_201 = _T_199 & ~reduced4CExtra; // @[MulAddRecFN.scala 137:44]
  assign _T_203 = mainAlignedSigC[2:0] != 3'h0; // @[MulAddRecFN.scala 138:39]
  assign _T_204 = _T_203 | reduced4CExtra; // @[MulAddRecFN.scala 138:44]
  assign _T_205 = doSubMags ? _T_201 : _T_204; // @[MulAddRecFN.scala 136:16]
  assign _T_206 = mainAlignedSigC[164:3]; // @[Cat.scala 30:58]
  assign alignedSigC = {_T_206,_T_205}; // @[Cat.scala 30:58]
  assign _T_210 = rawA_isNaN & ~rawA_sig[51]; // @[common.scala 81:46]
  assign _T_213 = rawB_isNaN & ~rawB_sig[51]; // @[common.scala 81:46]
  assign _T_214 = _T_210 | _T_213; // @[MulAddRecFN.scala 149:32]
  assign _T_217 = rawC_isNaN & ~rawC_sig[51]; // @[common.scala 81:46]
  assign _T_222 = $signed(sExpAlignedProd) - 14'sh35; // @[MulAddRecFN.scala 161:53]
  assign _T_223 = CIsDominant ? $signed({{1{rawC_sExp[12]}},rawC_sExp}) : $signed(_T_222); // @[MulAddRecFN.scala 161:12]
  assign io_mulAddA = rawA_sig[52:0]; // @[MulAddRecFN.scala 144:16]
  assign io_mulAddB = rawB_sig[52:0]; // @[MulAddRecFN.scala 145:16]
  assign io_mulAddC = alignedSigC[106:1]; // @[MulAddRecFN.scala 146:16]
  assign io_toPostMul_isSigNaNAny = _T_214 | _T_217; // @[MulAddRecFN.scala 148:30]
  assign io_toPostMul_isNaNAOrB = rawA_isNaN | rawB_isNaN; // @[MulAddRecFN.scala 151:28]
  assign io_toPostMul_isInfA = _T_16 & ~io_a[61]; // @[MulAddRecFN.scala 152:28]
  assign io_toPostMul_isZeroA = io_a[63:61] == 3'h0; // @[MulAddRecFN.scala 153:28]
  assign io_toPostMul_isInfB = _T_33 & ~io_b[61]; // @[MulAddRecFN.scala 154:28]
  assign io_toPostMul_isZeroB = io_b[63:61] == 3'h0; // @[MulAddRecFN.scala 155:28]
  assign io_toPostMul_signProd = _T_63 ^ io_op[1]; // @[MulAddRecFN.scala 156:28]
  assign io_toPostMul_isNaNC = _T_50 & io_c[61]; // @[MulAddRecFN.scala 157:28]
  assign io_toPostMul_isInfC = _T_50 & ~io_c[61]; // @[MulAddRecFN.scala 158:28]
  assign io_toPostMul_isZeroC = io_c[63:61] == 3'h0; // @[MulAddRecFN.scala 159:28]
  assign io_toPostMul_sExpSum = _T_223[12:0]; // @[MulAddRecFN.scala 160:28]
  assign io_toPostMul_doSubMags = _T_68 ^ io_op[0]; // @[MulAddRecFN.scala 162:28]
  assign io_toPostMul_CIsDominant = ~rawC_isZero & _T_76; // @[MulAddRecFN.scala 163:30]
  assign io_toPostMul_CDom_CAlignDist = CAlignDist[5:0]; // @[MulAddRecFN.scala 164:34]
  assign io_toPostMul_highAlignedSigC = alignedSigC[161:107]; // @[MulAddRecFN.scala 165:34]
  assign io_toPostMul_bit0AlignedSigC = alignedSigC[0]; // @[MulAddRecFN.scala 167:34]
  assign MulAddRecFNToRaw_preMul_1_covSum = 30'h0;
  assign io_covSum = MulAddRecFNToRaw_preMul_1_covSum;
  assign metaAssert = 1'h0;
endmodule
module MulAddRecFNToRaw_postMul_1(
  input          io_fromPreMul_isSigNaNAny,
  input          io_fromPreMul_isNaNAOrB,
  input          io_fromPreMul_isInfA,
  input          io_fromPreMul_isZeroA,
  input          io_fromPreMul_isInfB,
  input          io_fromPreMul_isZeroB,
  input          io_fromPreMul_signProd,
  input          io_fromPreMul_isNaNC,
  input          io_fromPreMul_isInfC,
  input          io_fromPreMul_isZeroC,
  input  [12:0]  io_fromPreMul_sExpSum,
  input          io_fromPreMul_doSubMags,
  input          io_fromPreMul_CIsDominant,
  input  [5:0]   io_fromPreMul_CDom_CAlignDist,
  input  [54:0]  io_fromPreMul_highAlignedSigC,
  input          io_fromPreMul_bit0AlignedSigC,
  input  [106:0] io_mulAddResult,
  input  [2:0]   io_roundingMode,
  output         io_invalidExc,
  output         io_rawOut_isNaN,
  output         io_rawOut_isInf,
  output         io_rawOut_isZero,
  output         io_rawOut_sign,
  output [12:0]  io_rawOut_sExp,
  output [55:0]  io_rawOut_sig,
  output [29:0]  io_covSum,
  output         metaAssert
);
  wire  roundingMode_min; // @[MulAddRecFN.scala 188:45]
  wire  CDom_sign; // @[MulAddRecFN.scala 192:42]
  wire [54:0] _T_11; // @[MulAddRecFN.scala 195:47]
  wire [54:0] _T_12; // @[MulAddRecFN.scala 194:16]
  wire [161:0] sigSum; // @[Cat.scala 30:58]
  wire [1:0] _T_15; // @[MulAddRecFN.scala 205:69]
  wire [12:0] _GEN_0; // @[MulAddRecFN.scala 205:43]
  wire [12:0] CDom_sExp; // @[MulAddRecFN.scala 205:43]
  wire [107:0] _T_23; // @[Cat.scala 30:58]
  wire [107:0] CDom_absSigSum; // @[MulAddRecFN.scala 207:12]
  wire  _T_26; // @[MulAddRecFN.scala 217:36]
  wire  _T_28; // @[MulAddRecFN.scala 218:37]
  wire  CDom_absSigSumExtra; // @[MulAddRecFN.scala 216:12]
  wire [170:0] _GEN_1; // @[MulAddRecFN.scala 221:24]
  wire [170:0] _T_29; // @[MulAddRecFN.scala 221:24]
  wire [57:0] CDom_mainSig; // @[MulAddRecFN.scala 221:56]
  wire [54:0] _T_31; // @[MulAddRecFN.scala 224:53]
  wire  _T_53; // @[primitives.scala 121:54]
  wire  _T_55; // @[primitives.scala 121:54]
  wire  _T_57; // @[primitives.scala 121:54]
  wire  _T_59; // @[primitives.scala 121:54]
  wire  _T_61; // @[primitives.scala 121:54]
  wire  _T_63; // @[primitives.scala 121:54]
  wire  _T_65; // @[primitives.scala 121:54]
  wire  _T_67; // @[primitives.scala 121:54]
  wire  _T_69; // @[primitives.scala 121:54]
  wire  _T_71; // @[primitives.scala 121:54]
  wire  _T_73; // @[primitives.scala 121:54]
  wire  _T_75; // @[primitives.scala 121:54]
  wire  _T_77; // @[primitives.scala 121:54]
  wire  _T_79; // @[primitives.scala 124:57]
  wire [6:0] _T_85; // @[primitives.scala 125:20]
  wire [13:0] _T_92; // @[primitives.scala 125:20]
  wire [16:0] _T_95; // @[primitives.scala 77:58]
  wire [7:0] _T_101; // @[Bitwise.scala 103:31]
  wire [7:0] _T_103; // @[Bitwise.scala 103:65]
  wire [7:0] _T_105; // @[Bitwise.scala 103:75]
  wire [7:0] _T_106; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_2; // @[Bitwise.scala 103:31]
  wire [7:0] _T_111; // @[Bitwise.scala 103:31]
  wire [7:0] _T_113; // @[Bitwise.scala 103:65]
  wire [7:0] _T_115; // @[Bitwise.scala 103:75]
  wire [7:0] _T_116; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_3; // @[Bitwise.scala 103:31]
  wire [7:0] _T_121; // @[Bitwise.scala 103:31]
  wire [7:0] _T_123; // @[Bitwise.scala 103:65]
  wire [7:0] _T_125; // @[Bitwise.scala 103:75]
  wire [7:0] _T_126; // @[Bitwise.scala 103:39]
  wire [12:0] _T_140; // @[Cat.scala 30:58]
  wire [13:0] _GEN_4; // @[MulAddRecFN.scala 224:72]
  wire [13:0] _T_141; // @[MulAddRecFN.scala 224:72]
  wire  CDom_reduced4SigExtra; // @[MulAddRecFN.scala 225:73]
  wire  _T_144; // @[MulAddRecFN.scala 228:32]
  wire  _T_145; // @[MulAddRecFN.scala 228:36]
  wire  _T_146; // @[MulAddRecFN.scala 228:61]
  wire [55:0] CDom_sig; // @[Cat.scala 30:58]
  wire  notCDom_signSigSum; // @[MulAddRecFN.scala 234:36]
  wire [108:0] _GEN_5; // @[MulAddRecFN.scala 238:41]
  wire [108:0] _T_151; // @[MulAddRecFN.scala 238:41]
  wire [108:0] notCDom_absSigSum; // @[MulAddRecFN.scala 236:12]
  wire  _T_214; // @[primitives.scala 104:54]
  wire  _T_216; // @[primitives.scala 104:54]
  wire  _T_218; // @[primitives.scala 104:54]
  wire  _T_220; // @[primitives.scala 104:54]
  wire  _T_222; // @[primitives.scala 104:54]
  wire  _T_224; // @[primitives.scala 104:54]
  wire  _T_226; // @[primitives.scala 104:54]
  wire  _T_228; // @[primitives.scala 104:54]
  wire  _T_230; // @[primitives.scala 104:54]
  wire  _T_232; // @[primitives.scala 104:54]
  wire  _T_234; // @[primitives.scala 104:54]
  wire  _T_236; // @[primitives.scala 104:54]
  wire  _T_238; // @[primitives.scala 104:54]
  wire  _T_240; // @[primitives.scala 104:54]
  wire  _T_242; // @[primitives.scala 104:54]
  wire  _T_244; // @[primitives.scala 104:54]
  wire  _T_246; // @[primitives.scala 104:54]
  wire  _T_248; // @[primitives.scala 104:54]
  wire  _T_250; // @[primitives.scala 104:54]
  wire  _T_252; // @[primitives.scala 104:54]
  wire  _T_254; // @[primitives.scala 104:54]
  wire  _T_256; // @[primitives.scala 104:54]
  wire  _T_258; // @[primitives.scala 104:54]
  wire  _T_260; // @[primitives.scala 104:54]
  wire  _T_262; // @[primitives.scala 104:54]
  wire  _T_264; // @[primitives.scala 104:54]
  wire  _T_266; // @[primitives.scala 104:54]
  wire  _T_268; // @[primitives.scala 104:54]
  wire  _T_270; // @[primitives.scala 104:54]
  wire  _T_272; // @[primitives.scala 104:54]
  wire  _T_274; // @[primitives.scala 104:54]
  wire  _T_276; // @[primitives.scala 104:54]
  wire  _T_278; // @[primitives.scala 104:54]
  wire  _T_280; // @[primitives.scala 104:54]
  wire  _T_282; // @[primitives.scala 104:54]
  wire  _T_284; // @[primitives.scala 104:54]
  wire  _T_286; // @[primitives.scala 104:54]
  wire  _T_288; // @[primitives.scala 104:54]
  wire  _T_290; // @[primitives.scala 104:54]
  wire  _T_292; // @[primitives.scala 104:54]
  wire  _T_294; // @[primitives.scala 104:54]
  wire  _T_296; // @[primitives.scala 104:54]
  wire  _T_298; // @[primitives.scala 104:54]
  wire  _T_300; // @[primitives.scala 104:54]
  wire  _T_302; // @[primitives.scala 104:54]
  wire  _T_304; // @[primitives.scala 104:54]
  wire  _T_306; // @[primitives.scala 104:54]
  wire  _T_308; // @[primitives.scala 104:54]
  wire  _T_310; // @[primitives.scala 104:54]
  wire  _T_312; // @[primitives.scala 104:54]
  wire  _T_314; // @[primitives.scala 104:54]
  wire  _T_316; // @[primitives.scala 104:54]
  wire  _T_318; // @[primitives.scala 104:54]
  wire  _T_320; // @[primitives.scala 104:54]
  wire [5:0] _T_327; // @[primitives.scala 108:20]
  wire [12:0] _T_334; // @[primitives.scala 108:20]
  wire [6:0] _T_340; // @[primitives.scala 108:20]
  wire [26:0] _T_348; // @[primitives.scala 108:20]
  wire [6:0] _T_354; // @[primitives.scala 108:20]
  wire [13:0] _T_361; // @[primitives.scala 108:20]
  wire [6:0] _T_367; // @[primitives.scala 108:20]
  wire [54:0] notCDom_reduced2AbsSigSum; // @[primitives.scala 108:20]
  wire [31:0] _T_380; // @[Bitwise.scala 103:31]
  wire [31:0] _T_382; // @[Bitwise.scala 103:65]
  wire [31:0] _T_384; // @[Bitwise.scala 103:75]
  wire [31:0] _T_385; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_6; // @[Bitwise.scala 103:31]
  wire [31:0] _T_390; // @[Bitwise.scala 103:31]
  wire [31:0] _T_392; // @[Bitwise.scala 103:65]
  wire [31:0] _T_394; // @[Bitwise.scala 103:75]
  wire [31:0] _T_395; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_7; // @[Bitwise.scala 103:31]
  wire [31:0] _T_400; // @[Bitwise.scala 103:31]
  wire [31:0] _T_402; // @[Bitwise.scala 103:65]
  wire [31:0] _T_404; // @[Bitwise.scala 103:75]
  wire [31:0] _T_405; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_8; // @[Bitwise.scala 103:31]
  wire [31:0] _T_410; // @[Bitwise.scala 103:31]
  wire [31:0] _T_412; // @[Bitwise.scala 103:65]
  wire [31:0] _T_414; // @[Bitwise.scala 103:75]
  wire [31:0] _T_415; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_9; // @[Bitwise.scala 103:31]
  wire [31:0] _T_420; // @[Bitwise.scala 103:31]
  wire [31:0] _T_422; // @[Bitwise.scala 103:65]
  wire [31:0] _T_424; // @[Bitwise.scala 103:75]
  wire [31:0] _T_425; // @[Bitwise.scala 103:39]
  wire [15:0] _T_431; // @[Bitwise.scala 103:31]
  wire [15:0] _T_433; // @[Bitwise.scala 103:65]
  wire [15:0] _T_435; // @[Bitwise.scala 103:75]
  wire [15:0] _T_436; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_10; // @[Bitwise.scala 103:31]
  wire [15:0] _T_441; // @[Bitwise.scala 103:31]
  wire [15:0] _T_443; // @[Bitwise.scala 103:65]
  wire [15:0] _T_445; // @[Bitwise.scala 103:75]
  wire [15:0] _T_446; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_11; // @[Bitwise.scala 103:31]
  wire [15:0] _T_451; // @[Bitwise.scala 103:31]
  wire [15:0] _T_453; // @[Bitwise.scala 103:65]
  wire [15:0] _T_455; // @[Bitwise.scala 103:75]
  wire [15:0] _T_456; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_12; // @[Bitwise.scala 103:31]
  wire [15:0] _T_461; // @[Bitwise.scala 103:31]
  wire [15:0] _T_463; // @[Bitwise.scala 103:65]
  wire [15:0] _T_465; // @[Bitwise.scala 103:75]
  wire [15:0] _T_466; // @[Bitwise.scala 103:39]
  wire [54:0] _T_487; // @[Cat.scala 30:58]
  wire [5:0] _T_543; // @[Mux.scala 31:69]
  wire [5:0] _T_544; // @[Mux.scala 31:69]
  wire [5:0] _T_545; // @[Mux.scala 31:69]
  wire [5:0] _T_546; // @[Mux.scala 31:69]
  wire [5:0] _T_547; // @[Mux.scala 31:69]
  wire [5:0] _T_548; // @[Mux.scala 31:69]
  wire [5:0] _T_549; // @[Mux.scala 31:69]
  wire [5:0] _T_550; // @[Mux.scala 31:69]
  wire [5:0] _T_551; // @[Mux.scala 31:69]
  wire [5:0] _T_552; // @[Mux.scala 31:69]
  wire [5:0] _T_553; // @[Mux.scala 31:69]
  wire [5:0] _T_554; // @[Mux.scala 31:69]
  wire [5:0] _T_555; // @[Mux.scala 31:69]
  wire [5:0] _T_556; // @[Mux.scala 31:69]
  wire [5:0] _T_557; // @[Mux.scala 31:69]
  wire [5:0] _T_558; // @[Mux.scala 31:69]
  wire [5:0] _T_559; // @[Mux.scala 31:69]
  wire [5:0] _T_560; // @[Mux.scala 31:69]
  wire [5:0] _T_561; // @[Mux.scala 31:69]
  wire [5:0] _T_562; // @[Mux.scala 31:69]
  wire [5:0] _T_563; // @[Mux.scala 31:69]
  wire [5:0] _T_564; // @[Mux.scala 31:69]
  wire [5:0] _T_565; // @[Mux.scala 31:69]
  wire [5:0] _T_566; // @[Mux.scala 31:69]
  wire [5:0] _T_567; // @[Mux.scala 31:69]
  wire [5:0] _T_568; // @[Mux.scala 31:69]
  wire [5:0] _T_569; // @[Mux.scala 31:69]
  wire [5:0] _T_570; // @[Mux.scala 31:69]
  wire [5:0] _T_571; // @[Mux.scala 31:69]
  wire [5:0] _T_572; // @[Mux.scala 31:69]
  wire [5:0] _T_573; // @[Mux.scala 31:69]
  wire [5:0] _T_574; // @[Mux.scala 31:69]
  wire [5:0] _T_575; // @[Mux.scala 31:69]
  wire [5:0] _T_576; // @[Mux.scala 31:69]
  wire [5:0] _T_577; // @[Mux.scala 31:69]
  wire [5:0] _T_578; // @[Mux.scala 31:69]
  wire [5:0] _T_579; // @[Mux.scala 31:69]
  wire [5:0] _T_580; // @[Mux.scala 31:69]
  wire [5:0] _T_581; // @[Mux.scala 31:69]
  wire [5:0] _T_582; // @[Mux.scala 31:69]
  wire [5:0] _T_583; // @[Mux.scala 31:69]
  wire [5:0] _T_584; // @[Mux.scala 31:69]
  wire [5:0] _T_585; // @[Mux.scala 31:69]
  wire [5:0] _T_586; // @[Mux.scala 31:69]
  wire [5:0] _T_587; // @[Mux.scala 31:69]
  wire [5:0] _T_588; // @[Mux.scala 31:69]
  wire [5:0] _T_589; // @[Mux.scala 31:69]
  wire [5:0] _T_590; // @[Mux.scala 31:69]
  wire [5:0] _T_591; // @[Mux.scala 31:69]
  wire [5:0] _T_592; // @[Mux.scala 31:69]
  wire [5:0] _T_593; // @[Mux.scala 31:69]
  wire [5:0] _T_594; // @[Mux.scala 31:69]
  wire [5:0] _T_595; // @[Mux.scala 31:69]
  wire [5:0] notCDom_normDistReduced2; // @[Mux.scala 31:69]
  wire [6:0] notCDom_nearNormDist; // @[MulAddRecFN.scala 242:56]
  wire [7:0] _T_596; // @[MulAddRecFN.scala 243:69]
  wire [12:0] _GEN_13; // @[MulAddRecFN.scala 243:46]
  wire [12:0] notCDom_sExp; // @[MulAddRecFN.scala 243:46]
  wire [235:0] _GEN_14; // @[MulAddRecFN.scala 245:27]
  wire [235:0] _T_599; // @[MulAddRecFN.scala 245:27]
  wire [57:0] notCDom_mainSig; // @[MulAddRecFN.scala 245:50]
  wire  _T_623; // @[primitives.scala 104:54]
  wire  _T_625; // @[primitives.scala 104:54]
  wire  _T_627; // @[primitives.scala 104:54]
  wire  _T_629; // @[primitives.scala 104:54]
  wire  _T_631; // @[primitives.scala 104:54]
  wire  _T_633; // @[primitives.scala 104:54]
  wire  _T_635; // @[primitives.scala 104:54]
  wire  _T_637; // @[primitives.scala 104:54]
  wire  _T_639; // @[primitives.scala 104:54]
  wire  _T_641; // @[primitives.scala 104:54]
  wire  _T_643; // @[primitives.scala 104:54]
  wire  _T_645; // @[primitives.scala 104:54]
  wire  _T_647; // @[primitives.scala 104:54]
  wire [6:0] _T_655; // @[primitives.scala 108:20]
  wire [13:0] _T_662; // @[primitives.scala 108:20]
  wire [32:0] _T_665; // @[primitives.scala 77:58]
  wire [7:0] _T_671; // @[Bitwise.scala 103:31]
  wire [7:0] _T_673; // @[Bitwise.scala 103:65]
  wire [7:0] _T_675; // @[Bitwise.scala 103:75]
  wire [7:0] _T_676; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_15; // @[Bitwise.scala 103:31]
  wire [7:0] _T_681; // @[Bitwise.scala 103:31]
  wire [7:0] _T_683; // @[Bitwise.scala 103:65]
  wire [7:0] _T_685; // @[Bitwise.scala 103:75]
  wire [7:0] _T_686; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_16; // @[Bitwise.scala 103:31]
  wire [7:0] _T_691; // @[Bitwise.scala 103:31]
  wire [7:0] _T_693; // @[Bitwise.scala 103:65]
  wire [7:0] _T_695; // @[Bitwise.scala 103:75]
  wire [7:0] _T_696; // @[Bitwise.scala 103:39]
  wire [12:0] _T_710; // @[Cat.scala 30:58]
  wire [13:0] _GEN_17; // @[MulAddRecFN.scala 249:78]
  wire [13:0] _T_711; // @[MulAddRecFN.scala 249:78]
  wire  notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 251:11]
  wire  _T_714; // @[MulAddRecFN.scala 254:35]
  wire  _T_715; // @[MulAddRecFN.scala 254:39]
  wire [55:0] notCDom_sig; // @[Cat.scala 30:58]
  wire  notCDom_completeCancellation; // @[MulAddRecFN.scala 257:50]
  wire  _T_717; // @[MulAddRecFN.scala 261:36]
  wire  notCDom_sign; // @[MulAddRecFN.scala 259:12]
  wire  notNaN_isInfProd; // @[MulAddRecFN.scala 266:49]
  wire  notNaN_isInfOut; // @[MulAddRecFN.scala 267:44]
  wire  _T_718; // @[MulAddRecFN.scala 269:32]
  wire  notNaN_addZeros; // @[MulAddRecFN.scala 269:58]
  wire  _T_719; // @[MulAddRecFN.scala 274:31]
  wire  _T_720; // @[MulAddRecFN.scala 273:35]
  wire  _T_721; // @[MulAddRecFN.scala 275:32]
  wire  _T_722; // @[MulAddRecFN.scala 274:57]
  wire  _T_725; // @[MulAddRecFN.scala 276:36]
  wire  _T_726; // @[MulAddRecFN.scala 277:61]
  wire  _T_727; // @[MulAddRecFN.scala 278:35]
  wire  _T_731; // @[MulAddRecFN.scala 285:42]
  wire  _T_733; // @[MulAddRecFN.scala 287:27]
  wire  _T_734; // @[MulAddRecFN.scala 288:31]
  wire  _T_735; // @[MulAddRecFN.scala 287:54]
  wire  _T_737; // @[MulAddRecFN.scala 289:26]
  wire  _T_738; // @[MulAddRecFN.scala 289:48]
  wire  _T_739; // @[MulAddRecFN.scala 290:36]
  wire  _T_740; // @[MulAddRecFN.scala 288:43]
  wire  _T_741; // @[MulAddRecFN.scala 291:26]
  wire  _T_742; // @[MulAddRecFN.scala 292:37]
  wire  _T_743; // @[MulAddRecFN.scala 291:46]
  wire  _T_744; // @[MulAddRecFN.scala 290:48]
  wire  _T_747; // @[MulAddRecFN.scala 293:28]
  wire  _T_748; // @[MulAddRecFN.scala 294:17]
  wire  _T_749; // @[MulAddRecFN.scala 293:49]
  wire [29:0] MulAddRecFNToRaw_postMul_1_covSum;
  assign roundingMode_min = io_roundingMode == 3'h2; // @[MulAddRecFN.scala 188:45]
  assign CDom_sign = io_fromPreMul_signProd ^ io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 192:42]
  assign _T_11 = io_fromPreMul_highAlignedSigC + 55'h1; // @[MulAddRecFN.scala 195:47]
  assign _T_12 = io_mulAddResult[106] ? _T_11 : io_fromPreMul_highAlignedSigC; // @[MulAddRecFN.scala 194:16]
  assign sigSum = {_T_12,io_mulAddResult[105:0],io_fromPreMul_bit0AlignedSigC}; // @[Cat.scala 30:58]
  assign _T_15 = {1'b0,$signed(io_fromPreMul_doSubMags)}; // @[MulAddRecFN.scala 205:69]
  assign _GEN_0 = {{11{_T_15[1]}},_T_15}; // @[MulAddRecFN.scala 205:43]
  assign CDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_0); // @[MulAddRecFN.scala 205:43]
  assign _T_23 = {1'h0,io_fromPreMul_highAlignedSigC[54:53],sigSum[159:55]}; // @[Cat.scala 30:58]
  assign CDom_absSigSum = io_fromPreMul_doSubMags ? ~sigSum[161:54] : _T_23; // @[MulAddRecFN.scala 207:12]
  assign _T_26 = ~sigSum[53:1] != 53'h0; // @[MulAddRecFN.scala 217:36]
  assign _T_28 = sigSum[54:1] != 54'h0; // @[MulAddRecFN.scala 218:37]
  assign CDom_absSigSumExtra = io_fromPreMul_doSubMags ? _T_26 : _T_28; // @[MulAddRecFN.scala 216:12]
  assign _GEN_1 = {{63'd0}, CDom_absSigSum}; // @[MulAddRecFN.scala 221:24]
  assign _T_29 = _GEN_1 << io_fromPreMul_CDom_CAlignDist; // @[MulAddRecFN.scala 221:24]
  assign CDom_mainSig = _T_29[107:50]; // @[MulAddRecFN.scala 221:56]
  assign _T_31 = {CDom_absSigSum[52:0], 2'h0}; // @[MulAddRecFN.scala 224:53]
  assign _T_53 = _T_31[3:0] != 4'h0; // @[primitives.scala 121:54]
  assign _T_55 = _T_31[7:4] != 4'h0; // @[primitives.scala 121:54]
  assign _T_57 = _T_31[11:8] != 4'h0; // @[primitives.scala 121:54]
  assign _T_59 = _T_31[15:12] != 4'h0; // @[primitives.scala 121:54]
  assign _T_61 = _T_31[19:16] != 4'h0; // @[primitives.scala 121:54]
  assign _T_63 = _T_31[23:20] != 4'h0; // @[primitives.scala 121:54]
  assign _T_65 = _T_31[27:24] != 4'h0; // @[primitives.scala 121:54]
  assign _T_67 = _T_31[31:28] != 4'h0; // @[primitives.scala 121:54]
  assign _T_69 = _T_31[35:32] != 4'h0; // @[primitives.scala 121:54]
  assign _T_71 = _T_31[39:36] != 4'h0; // @[primitives.scala 121:54]
  assign _T_73 = _T_31[43:40] != 4'h0; // @[primitives.scala 121:54]
  assign _T_75 = _T_31[47:44] != 4'h0; // @[primitives.scala 121:54]
  assign _T_77 = _T_31[51:48] != 4'h0; // @[primitives.scala 121:54]
  assign _T_79 = _T_31[54:52] != 3'h0; // @[primitives.scala 124:57]
  assign _T_85 = {_T_65,_T_63,_T_61,_T_59,_T_57,_T_55,_T_53}; // @[primitives.scala 125:20]
  assign _T_92 = {_T_79,_T_77,_T_75,_T_73,_T_71,_T_69,_T_67,_T_85}; // @[primitives.scala 125:20]
  assign _T_95 = -17'sh10000 >>> ~io_fromPreMul_CDom_CAlignDist[5:2]; // @[primitives.scala 77:58]
  assign _T_101 = {{4'd0}, _T_95[8:5]}; // @[Bitwise.scala 103:31]
  assign _T_103 = {_T_95[4:1], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_105 = _T_103 & 8'hf0; // @[Bitwise.scala 103:75]
  assign _T_106 = _T_101 | _T_105; // @[Bitwise.scala 103:39]
  assign _GEN_2 = {{2'd0}, _T_106[7:2]}; // @[Bitwise.scala 103:31]
  assign _T_111 = _GEN_2 & 8'h33; // @[Bitwise.scala 103:31]
  assign _T_113 = {_T_106[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_115 = _T_113 & 8'hcc; // @[Bitwise.scala 103:75]
  assign _T_116 = _T_111 | _T_115; // @[Bitwise.scala 103:39]
  assign _GEN_3 = {{1'd0}, _T_116[7:1]}; // @[Bitwise.scala 103:31]
  assign _T_121 = _GEN_3 & 8'h55; // @[Bitwise.scala 103:31]
  assign _T_123 = {_T_116[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_125 = _T_123 & 8'haa; // @[Bitwise.scala 103:75]
  assign _T_126 = _T_121 | _T_125; // @[Bitwise.scala 103:39]
  assign _T_140 = {_T_126,_T_95[9],_T_95[10],_T_95[11],_T_95[12],_T_95[13]}; // @[Cat.scala 30:58]
  assign _GEN_4 = {{1'd0}, _T_140}; // @[MulAddRecFN.scala 224:72]
  assign _T_141 = _T_92 & _GEN_4; // @[MulAddRecFN.scala 224:72]
  assign CDom_reduced4SigExtra = _T_141 != 14'h0; // @[MulAddRecFN.scala 225:73]
  assign _T_144 = CDom_mainSig[2:0] != 3'h0; // @[MulAddRecFN.scala 228:32]
  assign _T_145 = _T_144 | CDom_reduced4SigExtra; // @[MulAddRecFN.scala 228:36]
  assign _T_146 = _T_145 | CDom_absSigSumExtra; // @[MulAddRecFN.scala 228:61]
  assign CDom_sig = {CDom_mainSig[57:3],_T_146}; // @[Cat.scala 30:58]
  assign notCDom_signSigSum = sigSum[109]; // @[MulAddRecFN.scala 234:36]
  assign _GEN_5 = {{108'd0}, io_fromPreMul_doSubMags}; // @[MulAddRecFN.scala 238:41]
  assign _T_151 = sigSum[108:0] + _GEN_5; // @[MulAddRecFN.scala 238:41]
  assign notCDom_absSigSum = notCDom_signSigSum ? ~sigSum[108:0] : _T_151; // @[MulAddRecFN.scala 236:12]
  assign _T_214 = notCDom_absSigSum[1:0] != 2'h0; // @[primitives.scala 104:54]
  assign _T_216 = notCDom_absSigSum[3:2] != 2'h0; // @[primitives.scala 104:54]
  assign _T_218 = notCDom_absSigSum[5:4] != 2'h0; // @[primitives.scala 104:54]
  assign _T_220 = notCDom_absSigSum[7:6] != 2'h0; // @[primitives.scala 104:54]
  assign _T_222 = notCDom_absSigSum[9:8] != 2'h0; // @[primitives.scala 104:54]
  assign _T_224 = notCDom_absSigSum[11:10] != 2'h0; // @[primitives.scala 104:54]
  assign _T_226 = notCDom_absSigSum[13:12] != 2'h0; // @[primitives.scala 104:54]
  assign _T_228 = notCDom_absSigSum[15:14] != 2'h0; // @[primitives.scala 104:54]
  assign _T_230 = notCDom_absSigSum[17:16] != 2'h0; // @[primitives.scala 104:54]
  assign _T_232 = notCDom_absSigSum[19:18] != 2'h0; // @[primitives.scala 104:54]
  assign _T_234 = notCDom_absSigSum[21:20] != 2'h0; // @[primitives.scala 104:54]
  assign _T_236 = notCDom_absSigSum[23:22] != 2'h0; // @[primitives.scala 104:54]
  assign _T_238 = notCDom_absSigSum[25:24] != 2'h0; // @[primitives.scala 104:54]
  assign _T_240 = notCDom_absSigSum[27:26] != 2'h0; // @[primitives.scala 104:54]
  assign _T_242 = notCDom_absSigSum[29:28] != 2'h0; // @[primitives.scala 104:54]
  assign _T_244 = notCDom_absSigSum[31:30] != 2'h0; // @[primitives.scala 104:54]
  assign _T_246 = notCDom_absSigSum[33:32] != 2'h0; // @[primitives.scala 104:54]
  assign _T_248 = notCDom_absSigSum[35:34] != 2'h0; // @[primitives.scala 104:54]
  assign _T_250 = notCDom_absSigSum[37:36] != 2'h0; // @[primitives.scala 104:54]
  assign _T_252 = notCDom_absSigSum[39:38] != 2'h0; // @[primitives.scala 104:54]
  assign _T_254 = notCDom_absSigSum[41:40] != 2'h0; // @[primitives.scala 104:54]
  assign _T_256 = notCDom_absSigSum[43:42] != 2'h0; // @[primitives.scala 104:54]
  assign _T_258 = notCDom_absSigSum[45:44] != 2'h0; // @[primitives.scala 104:54]
  assign _T_260 = notCDom_absSigSum[47:46] != 2'h0; // @[primitives.scala 104:54]
  assign _T_262 = notCDom_absSigSum[49:48] != 2'h0; // @[primitives.scala 104:54]
  assign _T_264 = notCDom_absSigSum[51:50] != 2'h0; // @[primitives.scala 104:54]
  assign _T_266 = notCDom_absSigSum[53:52] != 2'h0; // @[primitives.scala 104:54]
  assign _T_268 = notCDom_absSigSum[55:54] != 2'h0; // @[primitives.scala 104:54]
  assign _T_270 = notCDom_absSigSum[57:56] != 2'h0; // @[primitives.scala 104:54]
  assign _T_272 = notCDom_absSigSum[59:58] != 2'h0; // @[primitives.scala 104:54]
  assign _T_274 = notCDom_absSigSum[61:60] != 2'h0; // @[primitives.scala 104:54]
  assign _T_276 = notCDom_absSigSum[63:62] != 2'h0; // @[primitives.scala 104:54]
  assign _T_278 = notCDom_absSigSum[65:64] != 2'h0; // @[primitives.scala 104:54]
  assign _T_280 = notCDom_absSigSum[67:66] != 2'h0; // @[primitives.scala 104:54]
  assign _T_282 = notCDom_absSigSum[69:68] != 2'h0; // @[primitives.scala 104:54]
  assign _T_284 = notCDom_absSigSum[71:70] != 2'h0; // @[primitives.scala 104:54]
  assign _T_286 = notCDom_absSigSum[73:72] != 2'h0; // @[primitives.scala 104:54]
  assign _T_288 = notCDom_absSigSum[75:74] != 2'h0; // @[primitives.scala 104:54]
  assign _T_290 = notCDom_absSigSum[77:76] != 2'h0; // @[primitives.scala 104:54]
  assign _T_292 = notCDom_absSigSum[79:78] != 2'h0; // @[primitives.scala 104:54]
  assign _T_294 = notCDom_absSigSum[81:80] != 2'h0; // @[primitives.scala 104:54]
  assign _T_296 = notCDom_absSigSum[83:82] != 2'h0; // @[primitives.scala 104:54]
  assign _T_298 = notCDom_absSigSum[85:84] != 2'h0; // @[primitives.scala 104:54]
  assign _T_300 = notCDom_absSigSum[87:86] != 2'h0; // @[primitives.scala 104:54]
  assign _T_302 = notCDom_absSigSum[89:88] != 2'h0; // @[primitives.scala 104:54]
  assign _T_304 = notCDom_absSigSum[91:90] != 2'h0; // @[primitives.scala 104:54]
  assign _T_306 = notCDom_absSigSum[93:92] != 2'h0; // @[primitives.scala 104:54]
  assign _T_308 = notCDom_absSigSum[95:94] != 2'h0; // @[primitives.scala 104:54]
  assign _T_310 = notCDom_absSigSum[97:96] != 2'h0; // @[primitives.scala 104:54]
  assign _T_312 = notCDom_absSigSum[99:98] != 2'h0; // @[primitives.scala 104:54]
  assign _T_314 = notCDom_absSigSum[101:100] != 2'h0; // @[primitives.scala 104:54]
  assign _T_316 = notCDom_absSigSum[103:102] != 2'h0; // @[primitives.scala 104:54]
  assign _T_318 = notCDom_absSigSum[105:104] != 2'h0; // @[primitives.scala 104:54]
  assign _T_320 = notCDom_absSigSum[107:106] != 2'h0; // @[primitives.scala 104:54]
  assign _T_327 = {_T_224,_T_222,_T_220,_T_218,_T_216,_T_214}; // @[primitives.scala 108:20]
  assign _T_334 = {_T_238,_T_236,_T_234,_T_232,_T_230,_T_228,_T_226,_T_327}; // @[primitives.scala 108:20]
  assign _T_340 = {_T_252,_T_250,_T_248,_T_246,_T_244,_T_242,_T_240}; // @[primitives.scala 108:20]
  assign _T_348 = {_T_266,_T_264,_T_262,_T_260,_T_258,_T_256,_T_254,_T_340,_T_334}; // @[primitives.scala 108:20]
  assign _T_354 = {_T_280,_T_278,_T_276,_T_274,_T_272,_T_270,_T_268}; // @[primitives.scala 108:20]
  assign _T_361 = {_T_294,_T_292,_T_290,_T_288,_T_286,_T_284,_T_282,_T_354}; // @[primitives.scala 108:20]
  assign _T_367 = {_T_308,_T_306,_T_304,_T_302,_T_300,_T_298,_T_296}; // @[primitives.scala 108:20]
  assign notCDom_reduced2AbsSigSum = {notCDom_absSigSum[108],_T_320,_T_318,_T_316,_T_314,_T_312,_T_310,_T_367,_T_361,_T_348}; // @[primitives.scala 108:20]
  assign _T_380 = {{16'd0}, notCDom_reduced2AbsSigSum[31:16]}; // @[Bitwise.scala 103:31]
  assign _T_382 = {notCDom_reduced2AbsSigSum[15:0], 16'h0}; // @[Bitwise.scala 103:65]
  assign _T_384 = _T_382 & 32'hffff0000; // @[Bitwise.scala 103:75]
  assign _T_385 = _T_380 | _T_384; // @[Bitwise.scala 103:39]
  assign _GEN_6 = {{8'd0}, _T_385[31:8]}; // @[Bitwise.scala 103:31]
  assign _T_390 = _GEN_6 & 32'hff00ff; // @[Bitwise.scala 103:31]
  assign _T_392 = {_T_385[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_394 = _T_392 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  assign _T_395 = _T_390 | _T_394; // @[Bitwise.scala 103:39]
  assign _GEN_7 = {{4'd0}, _T_395[31:4]}; // @[Bitwise.scala 103:31]
  assign _T_400 = _GEN_7 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  assign _T_402 = {_T_395[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_404 = _T_402 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  assign _T_405 = _T_400 | _T_404; // @[Bitwise.scala 103:39]
  assign _GEN_8 = {{2'd0}, _T_405[31:2]}; // @[Bitwise.scala 103:31]
  assign _T_410 = _GEN_8 & 32'h33333333; // @[Bitwise.scala 103:31]
  assign _T_412 = {_T_405[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_414 = _T_412 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  assign _T_415 = _T_410 | _T_414; // @[Bitwise.scala 103:39]
  assign _GEN_9 = {{1'd0}, _T_415[31:1]}; // @[Bitwise.scala 103:31]
  assign _T_420 = _GEN_9 & 32'h55555555; // @[Bitwise.scala 103:31]
  assign _T_422 = {_T_415[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_424 = _T_422 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  assign _T_425 = _T_420 | _T_424; // @[Bitwise.scala 103:39]
  assign _T_431 = {{8'd0}, notCDom_reduced2AbsSigSum[47:40]}; // @[Bitwise.scala 103:31]
  assign _T_433 = {notCDom_reduced2AbsSigSum[39:32], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_435 = _T_433 & 16'hff00; // @[Bitwise.scala 103:75]
  assign _T_436 = _T_431 | _T_435; // @[Bitwise.scala 103:39]
  assign _GEN_10 = {{4'd0}, _T_436[15:4]}; // @[Bitwise.scala 103:31]
  assign _T_441 = _GEN_10 & 16'hf0f; // @[Bitwise.scala 103:31]
  assign _T_443 = {_T_436[11:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_445 = _T_443 & 16'hf0f0; // @[Bitwise.scala 103:75]
  assign _T_446 = _T_441 | _T_445; // @[Bitwise.scala 103:39]
  assign _GEN_11 = {{2'd0}, _T_446[15:2]}; // @[Bitwise.scala 103:31]
  assign _T_451 = _GEN_11 & 16'h3333; // @[Bitwise.scala 103:31]
  assign _T_453 = {_T_446[13:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_455 = _T_453 & 16'hcccc; // @[Bitwise.scala 103:75]
  assign _T_456 = _T_451 | _T_455; // @[Bitwise.scala 103:39]
  assign _GEN_12 = {{1'd0}, _T_456[15:1]}; // @[Bitwise.scala 103:31]
  assign _T_461 = _GEN_12 & 16'h5555; // @[Bitwise.scala 103:31]
  assign _T_463 = {_T_456[14:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_465 = _T_463 & 16'haaaa; // @[Bitwise.scala 103:75]
  assign _T_466 = _T_461 | _T_465; // @[Bitwise.scala 103:39]
  assign _T_487 = {_T_425,_T_466,notCDom_reduced2AbsSigSum[48],notCDom_reduced2AbsSigSum[49],notCDom_reduced2AbsSigSum[50],notCDom_reduced2AbsSigSum[51],notCDom_reduced2AbsSigSum[52],notCDom_reduced2AbsSigSum[53],notCDom_reduced2AbsSigSum[54]}; // @[Cat.scala 30:58]
  assign _T_543 = _T_487[53] ? 6'h35 : 6'h36; // @[Mux.scala 31:69]
  assign _T_544 = _T_487[52] ? 6'h34 : _T_543; // @[Mux.scala 31:69]
  assign _T_545 = _T_487[51] ? 6'h33 : _T_544; // @[Mux.scala 31:69]
  assign _T_546 = _T_487[50] ? 6'h32 : _T_545; // @[Mux.scala 31:69]
  assign _T_547 = _T_487[49] ? 6'h31 : _T_546; // @[Mux.scala 31:69]
  assign _T_548 = _T_487[48] ? 6'h30 : _T_547; // @[Mux.scala 31:69]
  assign _T_549 = _T_487[47] ? 6'h2f : _T_548; // @[Mux.scala 31:69]
  assign _T_550 = _T_487[46] ? 6'h2e : _T_549; // @[Mux.scala 31:69]
  assign _T_551 = _T_487[45] ? 6'h2d : _T_550; // @[Mux.scala 31:69]
  assign _T_552 = _T_487[44] ? 6'h2c : _T_551; // @[Mux.scala 31:69]
  assign _T_553 = _T_487[43] ? 6'h2b : _T_552; // @[Mux.scala 31:69]
  assign _T_554 = _T_487[42] ? 6'h2a : _T_553; // @[Mux.scala 31:69]
  assign _T_555 = _T_487[41] ? 6'h29 : _T_554; // @[Mux.scala 31:69]
  assign _T_556 = _T_487[40] ? 6'h28 : _T_555; // @[Mux.scala 31:69]
  assign _T_557 = _T_487[39] ? 6'h27 : _T_556; // @[Mux.scala 31:69]
  assign _T_558 = _T_487[38] ? 6'h26 : _T_557; // @[Mux.scala 31:69]
  assign _T_559 = _T_487[37] ? 6'h25 : _T_558; // @[Mux.scala 31:69]
  assign _T_560 = _T_487[36] ? 6'h24 : _T_559; // @[Mux.scala 31:69]
  assign _T_561 = _T_487[35] ? 6'h23 : _T_560; // @[Mux.scala 31:69]
  assign _T_562 = _T_487[34] ? 6'h22 : _T_561; // @[Mux.scala 31:69]
  assign _T_563 = _T_487[33] ? 6'h21 : _T_562; // @[Mux.scala 31:69]
  assign _T_564 = _T_487[32] ? 6'h20 : _T_563; // @[Mux.scala 31:69]
  assign _T_565 = _T_487[31] ? 6'h1f : _T_564; // @[Mux.scala 31:69]
  assign _T_566 = _T_487[30] ? 6'h1e : _T_565; // @[Mux.scala 31:69]
  assign _T_567 = _T_487[29] ? 6'h1d : _T_566; // @[Mux.scala 31:69]
  assign _T_568 = _T_487[28] ? 6'h1c : _T_567; // @[Mux.scala 31:69]
  assign _T_569 = _T_487[27] ? 6'h1b : _T_568; // @[Mux.scala 31:69]
  assign _T_570 = _T_487[26] ? 6'h1a : _T_569; // @[Mux.scala 31:69]
  assign _T_571 = _T_487[25] ? 6'h19 : _T_570; // @[Mux.scala 31:69]
  assign _T_572 = _T_487[24] ? 6'h18 : _T_571; // @[Mux.scala 31:69]
  assign _T_573 = _T_487[23] ? 6'h17 : _T_572; // @[Mux.scala 31:69]
  assign _T_574 = _T_487[22] ? 6'h16 : _T_573; // @[Mux.scala 31:69]
  assign _T_575 = _T_487[21] ? 6'h15 : _T_574; // @[Mux.scala 31:69]
  assign _T_576 = _T_487[20] ? 6'h14 : _T_575; // @[Mux.scala 31:69]
  assign _T_577 = _T_487[19] ? 6'h13 : _T_576; // @[Mux.scala 31:69]
  assign _T_578 = _T_487[18] ? 6'h12 : _T_577; // @[Mux.scala 31:69]
  assign _T_579 = _T_487[17] ? 6'h11 : _T_578; // @[Mux.scala 31:69]
  assign _T_580 = _T_487[16] ? 6'h10 : _T_579; // @[Mux.scala 31:69]
  assign _T_581 = _T_487[15] ? 6'hf : _T_580; // @[Mux.scala 31:69]
  assign _T_582 = _T_487[14] ? 6'he : _T_581; // @[Mux.scala 31:69]
  assign _T_583 = _T_487[13] ? 6'hd : _T_582; // @[Mux.scala 31:69]
  assign _T_584 = _T_487[12] ? 6'hc : _T_583; // @[Mux.scala 31:69]
  assign _T_585 = _T_487[11] ? 6'hb : _T_584; // @[Mux.scala 31:69]
  assign _T_586 = _T_487[10] ? 6'ha : _T_585; // @[Mux.scala 31:69]
  assign _T_587 = _T_487[9] ? 6'h9 : _T_586; // @[Mux.scala 31:69]
  assign _T_588 = _T_487[8] ? 6'h8 : _T_587; // @[Mux.scala 31:69]
  assign _T_589 = _T_487[7] ? 6'h7 : _T_588; // @[Mux.scala 31:69]
  assign _T_590 = _T_487[6] ? 6'h6 : _T_589; // @[Mux.scala 31:69]
  assign _T_591 = _T_487[5] ? 6'h5 : _T_590; // @[Mux.scala 31:69]
  assign _T_592 = _T_487[4] ? 6'h4 : _T_591; // @[Mux.scala 31:69]
  assign _T_593 = _T_487[3] ? 6'h3 : _T_592; // @[Mux.scala 31:69]
  assign _T_594 = _T_487[2] ? 6'h2 : _T_593; // @[Mux.scala 31:69]
  assign _T_595 = _T_487[1] ? 6'h1 : _T_594; // @[Mux.scala 31:69]
  assign notCDom_normDistReduced2 = _T_487[0] ? 6'h0 : _T_595; // @[Mux.scala 31:69]
  assign notCDom_nearNormDist = {notCDom_normDistReduced2, 1'h0}; // @[MulAddRecFN.scala 242:56]
  assign _T_596 = {1'b0,$signed(notCDom_nearNormDist)}; // @[MulAddRecFN.scala 243:69]
  assign _GEN_13 = {{5{_T_596[7]}},_T_596}; // @[MulAddRecFN.scala 243:46]
  assign notCDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_13); // @[MulAddRecFN.scala 243:46]
  assign _GEN_14 = {{127'd0}, notCDom_absSigSum}; // @[MulAddRecFN.scala 245:27]
  assign _T_599 = _GEN_14 << notCDom_nearNormDist; // @[MulAddRecFN.scala 245:27]
  assign notCDom_mainSig = _T_599[109:52]; // @[MulAddRecFN.scala 245:50]
  assign _T_623 = notCDom_reduced2AbsSigSum[1:0] != 2'h0; // @[primitives.scala 104:54]
  assign _T_625 = notCDom_reduced2AbsSigSum[3:2] != 2'h0; // @[primitives.scala 104:54]
  assign _T_627 = notCDom_reduced2AbsSigSum[5:4] != 2'h0; // @[primitives.scala 104:54]
  assign _T_629 = notCDom_reduced2AbsSigSum[7:6] != 2'h0; // @[primitives.scala 104:54]
  assign _T_631 = notCDom_reduced2AbsSigSum[9:8] != 2'h0; // @[primitives.scala 104:54]
  assign _T_633 = notCDom_reduced2AbsSigSum[11:10] != 2'h0; // @[primitives.scala 104:54]
  assign _T_635 = notCDom_reduced2AbsSigSum[13:12] != 2'h0; // @[primitives.scala 104:54]
  assign _T_637 = notCDom_reduced2AbsSigSum[15:14] != 2'h0; // @[primitives.scala 104:54]
  assign _T_639 = notCDom_reduced2AbsSigSum[17:16] != 2'h0; // @[primitives.scala 104:54]
  assign _T_641 = notCDom_reduced2AbsSigSum[19:18] != 2'h0; // @[primitives.scala 104:54]
  assign _T_643 = notCDom_reduced2AbsSigSum[21:20] != 2'h0; // @[primitives.scala 104:54]
  assign _T_645 = notCDom_reduced2AbsSigSum[23:22] != 2'h0; // @[primitives.scala 104:54]
  assign _T_647 = notCDom_reduced2AbsSigSum[25:24] != 2'h0; // @[primitives.scala 104:54]
  assign _T_655 = {_T_635,_T_633,_T_631,_T_629,_T_627,_T_625,_T_623}; // @[primitives.scala 108:20]
  assign _T_662 = {notCDom_reduced2AbsSigSum[26],_T_647,_T_645,_T_643,_T_641,_T_639,_T_637,_T_655}; // @[primitives.scala 108:20]
  assign _T_665 = -33'sh100000000 >>> ~notCDom_normDistReduced2[5:1]; // @[primitives.scala 77:58]
  assign _T_671 = {{4'd0}, _T_665[8:5]}; // @[Bitwise.scala 103:31]
  assign _T_673 = {_T_665[4:1], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_675 = _T_673 & 8'hf0; // @[Bitwise.scala 103:75]
  assign _T_676 = _T_671 | _T_675; // @[Bitwise.scala 103:39]
  assign _GEN_15 = {{2'd0}, _T_676[7:2]}; // @[Bitwise.scala 103:31]
  assign _T_681 = _GEN_15 & 8'h33; // @[Bitwise.scala 103:31]
  assign _T_683 = {_T_676[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_685 = _T_683 & 8'hcc; // @[Bitwise.scala 103:75]
  assign _T_686 = _T_681 | _T_685; // @[Bitwise.scala 103:39]
  assign _GEN_16 = {{1'd0}, _T_686[7:1]}; // @[Bitwise.scala 103:31]
  assign _T_691 = _GEN_16 & 8'h55; // @[Bitwise.scala 103:31]
  assign _T_693 = {_T_686[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_695 = _T_693 & 8'haa; // @[Bitwise.scala 103:75]
  assign _T_696 = _T_691 | _T_695; // @[Bitwise.scala 103:39]
  assign _T_710 = {_T_696,_T_665[9],_T_665[10],_T_665[11],_T_665[12],_T_665[13]}; // @[Cat.scala 30:58]
  assign _GEN_17 = {{1'd0}, _T_710}; // @[MulAddRecFN.scala 249:78]
  assign _T_711 = _T_662 & _GEN_17; // @[MulAddRecFN.scala 249:78]
  assign notCDom_reduced4SigExtra = _T_711 != 14'h0; // @[MulAddRecFN.scala 251:11]
  assign _T_714 = notCDom_mainSig[2:0] != 3'h0; // @[MulAddRecFN.scala 254:35]
  assign _T_715 = _T_714 | notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 254:39]
  assign notCDom_sig = {notCDom_mainSig[57:3],_T_715}; // @[Cat.scala 30:58]
  assign notCDom_completeCancellation = notCDom_sig[55:54] == 2'h0; // @[MulAddRecFN.scala 257:50]
  assign _T_717 = io_fromPreMul_signProd ^ notCDom_signSigSum; // @[MulAddRecFN.scala 261:36]
  assign notCDom_sign = notCDom_completeCancellation ? roundingMode_min : _T_717; // @[MulAddRecFN.scala 259:12]
  assign notNaN_isInfProd = io_fromPreMul_isInfA | io_fromPreMul_isInfB; // @[MulAddRecFN.scala 266:49]
  assign notNaN_isInfOut = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 267:44]
  assign _T_718 = io_fromPreMul_isZeroA | io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 269:32]
  assign notNaN_addZeros = _T_718 & io_fromPreMul_isZeroC; // @[MulAddRecFN.scala 269:58]
  assign _T_719 = io_fromPreMul_isInfA & io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 274:31]
  assign _T_720 = io_fromPreMul_isSigNaNAny | _T_719; // @[MulAddRecFN.scala 273:35]
  assign _T_721 = io_fromPreMul_isZeroA & io_fromPreMul_isInfB; // @[MulAddRecFN.scala 275:32]
  assign _T_722 = _T_720 | _T_721; // @[MulAddRecFN.scala 274:57]
  assign _T_725 = ~io_fromPreMul_isNaNAOrB & notNaN_isInfProd; // @[MulAddRecFN.scala 276:36]
  assign _T_726 = _T_725 & io_fromPreMul_isInfC; // @[MulAddRecFN.scala 277:61]
  assign _T_727 = _T_726 & io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 278:35]
  assign _T_731 = ~io_fromPreMul_CIsDominant & notCDom_completeCancellation; // @[MulAddRecFN.scala 285:42]
  assign _T_733 = notNaN_isInfProd & io_fromPreMul_signProd; // @[MulAddRecFN.scala 287:27]
  assign _T_734 = io_fromPreMul_isInfC & CDom_sign; // @[MulAddRecFN.scala 288:31]
  assign _T_735 = _T_733 | _T_734; // @[MulAddRecFN.scala 287:54]
  assign _T_737 = notNaN_addZeros & ~roundingMode_min; // @[MulAddRecFN.scala 289:26]
  assign _T_738 = _T_737 & io_fromPreMul_signProd; // @[MulAddRecFN.scala 289:48]
  assign _T_739 = _T_738 & CDom_sign; // @[MulAddRecFN.scala 290:36]
  assign _T_740 = _T_735 | _T_739; // @[MulAddRecFN.scala 288:43]
  assign _T_741 = notNaN_addZeros & roundingMode_min; // @[MulAddRecFN.scala 291:26]
  assign _T_742 = io_fromPreMul_signProd | CDom_sign; // @[MulAddRecFN.scala 292:37]
  assign _T_743 = _T_741 & _T_742; // @[MulAddRecFN.scala 291:46]
  assign _T_744 = _T_740 | _T_743; // @[MulAddRecFN.scala 290:48]
  assign _T_747 = ~notNaN_isInfOut & ~notNaN_addZeros; // @[MulAddRecFN.scala 293:28]
  assign _T_748 = io_fromPreMul_CIsDominant ? CDom_sign : notCDom_sign; // @[MulAddRecFN.scala 294:17]
  assign _T_749 = _T_747 & _T_748; // @[MulAddRecFN.scala 293:49]
  assign io_invalidExc = _T_722 | _T_727; // @[MulAddRecFN.scala 272:19]
  assign io_rawOut_isNaN = io_fromPreMul_isNaNAOrB | io_fromPreMul_isNaNC; // @[MulAddRecFN.scala 280:21]
  assign io_rawOut_isInf = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 281:21]
  assign io_rawOut_isZero = notNaN_addZeros | _T_731; // @[MulAddRecFN.scala 283:22]
  assign io_rawOut_sign = _T_744 | _T_749; // @[MulAddRecFN.scala 286:20]
  assign io_rawOut_sExp = io_fromPreMul_CIsDominant ? $signed(CDom_sExp) : $signed(notCDom_sExp); // @[MulAddRecFN.scala 295:20]
  assign io_rawOut_sig = io_fromPreMul_CIsDominant ? CDom_sig : notCDom_sig; // @[MulAddRecFN.scala 296:19]
  assign MulAddRecFNToRaw_postMul_1_covSum = 30'h0;
  assign io_covSum = MulAddRecFNToRaw_postMul_1_covSum;
  assign metaAssert = 1'h0;
endmodule
module RoundAnyRawFNToRecFN_5(
  input         io_invalidExc,
  input         io_infiniteExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [9:0]  io_in_sExp,
  input  [26:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire  _T_11; // @[RoundAnyRawFNToRecFN.scala 96:27]
  wire  _T_13; // @[RoundAnyRawFNToRecFN.scala 96:63]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42]
  wire  doShiftSigDown1; // @[RoundAnyRawFNToRecFN.scala 118:61]
  wire  _T_22; // @[primitives.scala 57:25]
  wire  _T_24; // @[primitives.scala 57:25]
  wire  _T_26; // @[primitives.scala 57:25]
  wire [5:0] _T_27; // @[primitives.scala 58:26]
  wire [64:0] _T_28; // @[primitives.scala 77:58]
  wire [15:0] _T_34; // @[Bitwise.scala 103:31]
  wire [15:0] _T_36; // @[Bitwise.scala 103:65]
  wire [15:0] _T_38; // @[Bitwise.scala 103:75]
  wire [15:0] _T_39; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_0; // @[Bitwise.scala 103:31]
  wire [15:0] _T_44; // @[Bitwise.scala 103:31]
  wire [15:0] _T_46; // @[Bitwise.scala 103:65]
  wire [15:0] _T_48; // @[Bitwise.scala 103:75]
  wire [15:0] _T_49; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_1; // @[Bitwise.scala 103:31]
  wire [15:0] _T_54; // @[Bitwise.scala 103:31]
  wire [15:0] _T_56; // @[Bitwise.scala 103:65]
  wire [15:0] _T_58; // @[Bitwise.scala 103:75]
  wire [15:0] _T_59; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_2; // @[Bitwise.scala 103:31]
  wire [15:0] _T_64; // @[Bitwise.scala 103:31]
  wire [15:0] _T_66; // @[Bitwise.scala 103:65]
  wire [15:0] _T_68; // @[Bitwise.scala 103:75]
  wire [15:0] _T_69; // @[Bitwise.scala 103:39]
  wire [21:0] _T_86; // @[Cat.scala 30:58]
  wire [21:0] _T_88; // @[primitives.scala 74:21]
  wire [24:0] _T_90; // @[Cat.scala 30:58]
  wire [2:0] _T_100; // @[Cat.scala 30:58]
  wire [2:0] _T_101; // @[primitives.scala 61:24]
  wire [24:0] _T_102; // @[primitives.scala 66:24]
  wire [24:0] _T_103; // @[primitives.scala 61:24]
  wire [24:0] _GEN_3; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [24:0] _T_104; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [26:0] _T_105; // @[Cat.scala 30:58]
  wire [26:0] _T_107; // @[Cat.scala 30:58]
  wire [26:0] _T_109; // @[RoundAnyRawFNToRecFN.scala 161:46]
  wire [26:0] _T_110; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  _T_111; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [26:0] _T_112; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  _T_113; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  _T_114; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire  _T_115; // @[RoundAnyRawFNToRecFN.scala 167:38]
  wire  _T_116; // @[RoundAnyRawFNToRecFN.scala 167:67]
  wire  _T_117; // @[RoundAnyRawFNToRecFN.scala 169:29]
  wire  _T_118; // @[RoundAnyRawFNToRecFN.scala 168:31]
  wire [26:0] _T_119; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [25:0] _T_121; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _T_122; // @[RoundAnyRawFNToRecFN.scala 173:49]
  wire  _T_124; // @[RoundAnyRawFNToRecFN.scala 173:64]
  wire [25:0] _T_126; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [25:0] _T_128; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [26:0] _T_130; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire  _T_132; // @[RoundAnyRawFNToRecFN.scala 179:42]
  wire [25:0] _T_134; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [25:0] _GEN_4; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] _T_135; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] _T_136; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _T_138; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [9:0] _GEN_5; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [10:0] _T_139; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [8:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [22:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 187:16]
  wire [3:0] _T_144; // @[RoundAnyRawFNToRecFN.scala 194:30]
  wire  common_overflow; // @[RoundAnyRawFNToRecFN.scala 194:50]
  wire  common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 198:31]
  wire  _T_149; // @[RoundAnyRawFNToRecFN.scala 201:16]
  wire  _T_151; // @[RoundAnyRawFNToRecFN.scala 203:30]
  wire  _T_153; // @[RoundAnyRawFNToRecFN.scala 203:70]
  wire  _T_154; // @[RoundAnyRawFNToRecFN.scala 203:49]
  wire  _T_156; // @[RoundAnyRawFNToRecFN.scala 205:67]
  wire  _T_157; // @[RoundAnyRawFNToRecFN.scala 207:29]
  wire  _T_158; // @[RoundAnyRawFNToRecFN.scala 206:46]
  wire  _T_161; // @[RoundAnyRawFNToRecFN.scala 209:16]
  wire [1:0] _T_162; // @[RoundAnyRawFNToRecFN.scala 218:48]
  wire  _T_163; // @[RoundAnyRawFNToRecFN.scala 218:62]
  wire  _T_164; // @[RoundAnyRawFNToRecFN.scala 218:32]
  wire  _T_167; // @[RoundAnyRawFNToRecFN.scala 219:30]
  wire  _T_168; // @[RoundAnyRawFNToRecFN.scala 218:74]
  wire  _T_172; // @[RoundAnyRawFNToRecFN.scala 221:39]
  wire  _T_174; // @[RoundAnyRawFNToRecFN.scala 220:77]
  wire  _T_175; // @[RoundAnyRawFNToRecFN.scala 224:38]
  wire  _T_176; // @[RoundAnyRawFNToRecFN.scala 225:45]
  wire  _T_177; // @[RoundAnyRawFNToRecFN.scala 225:60]
  wire  _T_179; // @[RoundAnyRawFNToRecFN.scala 219:76]
  wire  common_underflow; // @[RoundAnyRawFNToRecFN.scala 215:40]
  wire  common_inexact; // @[RoundAnyRawFNToRecFN.scala 228:49]
  wire  isNaNOut; // @[RoundAnyRawFNToRecFN.scala 233:34]
  wire  notNaN_isSpecialInfOut; // @[RoundAnyRawFNToRecFN.scala 234:49]
  wire  _T_184; // @[RoundAnyRawFNToRecFN.scala 235:33]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:61]
  wire  overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  wire  underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  wire  _T_186; // @[RoundAnyRawFNToRecFN.scala 238:43]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:28]
  wire  overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  wire  _T_188; // @[RoundAnyRawFNToRecFN.scala 243:20]
  wire  _T_189; // @[RoundAnyRawFNToRecFN.scala 243:60]
  wire  pegMinNonzeroMagOut; // @[RoundAnyRawFNToRecFN.scala 243:45]
  wire  pegMaxFiniteMagOut; // @[RoundAnyRawFNToRecFN.scala 244:39]
  wire  _T_191; // @[RoundAnyRawFNToRecFN.scala 246:45]
  wire  notNaN_isInfOut; // @[RoundAnyRawFNToRecFN.scala 246:32]
  wire  signOut; // @[RoundAnyRawFNToRecFN.scala 248:22]
  wire  _T_192; // @[RoundAnyRawFNToRecFN.scala 251:32]
  wire [8:0] _T_193; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [8:0] _T_195; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [8:0] _T_197; // @[RoundAnyRawFNToRecFN.scala 255:18]
  wire [8:0] _T_199; // @[RoundAnyRawFNToRecFN.scala 254:17]
  wire [8:0] _T_200; // @[RoundAnyRawFNToRecFN.scala 259:18]
  wire [8:0] _T_202; // @[RoundAnyRawFNToRecFN.scala 258:17]
  wire [8:0] _T_203; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [8:0] _T_205; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [8:0] _T_206; // @[RoundAnyRawFNToRecFN.scala 267:16]
  wire [8:0] _T_207; // @[RoundAnyRawFNToRecFN.scala 266:18]
  wire [8:0] _T_208; // @[RoundAnyRawFNToRecFN.scala 271:16]
  wire [8:0] _T_209; // @[RoundAnyRawFNToRecFN.scala 270:15]
  wire [8:0] _T_210; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [8:0] _T_211; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [8:0] _T_212; // @[RoundAnyRawFNToRecFN.scala 276:16]
  wire [8:0] expOut; // @[RoundAnyRawFNToRecFN.scala 275:77]
  wire  _T_213; // @[RoundAnyRawFNToRecFN.scala 278:22]
  wire  _T_214; // @[RoundAnyRawFNToRecFN.scala 278:38]
  wire [22:0] _T_215; // @[RoundAnyRawFNToRecFN.scala 279:16]
  wire [22:0] _T_216; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [22:0] _T_218; // @[Bitwise.scala 72:12]
  wire [22:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 281:11]
  wire [9:0] _T_219; // @[Cat.scala 30:58]
  wire [1:0] _T_221; // @[Cat.scala 30:58]
  wire [2:0] _T_223; // @[Cat.scala 30:58]
  wire [29:0] RoundAnyRawFNToRecFN_5_covSum;
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53]
  assign roundingMode_odd = io_roundingMode == 3'h5; // @[RoundAnyRawFNToRecFN.scala 93:53]
  assign _T_11 = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27]
  assign _T_13 = roundingMode_max & ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:63]
  assign roundMagUp = _T_11 | _T_13; // @[RoundAnyRawFNToRecFN.scala 96:42]
  assign doShiftSigDown1 = io_in_sig[26]; // @[RoundAnyRawFNToRecFN.scala 118:61]
  assign _T_22 = ~io_in_sExp[8]; // @[primitives.scala 57:25]
  assign _T_24 = ~io_in_sExp[7]; // @[primitives.scala 57:25]
  assign _T_26 = ~io_in_sExp[6]; // @[primitives.scala 57:25]
  assign _T_27 = ~io_in_sExp[5:0]; // @[primitives.scala 58:26]
  assign _T_28 = -65'sh10000000000000000 >>> _T_27; // @[primitives.scala 77:58]
  assign _T_34 = {{8'd0}, _T_28[57:50]}; // @[Bitwise.scala 103:31]
  assign _T_36 = {_T_28[49:42], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_38 = _T_36 & 16'hff00; // @[Bitwise.scala 103:75]
  assign _T_39 = _T_34 | _T_38; // @[Bitwise.scala 103:39]
  assign _GEN_0 = {{4'd0}, _T_39[15:4]}; // @[Bitwise.scala 103:31]
  assign _T_44 = _GEN_0 & 16'hf0f; // @[Bitwise.scala 103:31]
  assign _T_46 = {_T_39[11:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_48 = _T_46 & 16'hf0f0; // @[Bitwise.scala 103:75]
  assign _T_49 = _T_44 | _T_48; // @[Bitwise.scala 103:39]
  assign _GEN_1 = {{2'd0}, _T_49[15:2]}; // @[Bitwise.scala 103:31]
  assign _T_54 = _GEN_1 & 16'h3333; // @[Bitwise.scala 103:31]
  assign _T_56 = {_T_49[13:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_58 = _T_56 & 16'hcccc; // @[Bitwise.scala 103:75]
  assign _T_59 = _T_54 | _T_58; // @[Bitwise.scala 103:39]
  assign _GEN_2 = {{1'd0}, _T_59[15:1]}; // @[Bitwise.scala 103:31]
  assign _T_64 = _GEN_2 & 16'h5555; // @[Bitwise.scala 103:31]
  assign _T_66 = {_T_59[14:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_68 = _T_66 & 16'haaaa; // @[Bitwise.scala 103:75]
  assign _T_69 = _T_64 | _T_68; // @[Bitwise.scala 103:39]
  assign _T_86 = {_T_69,_T_28[58],_T_28[59],_T_28[60],_T_28[61],_T_28[62],_T_28[63]}; // @[Cat.scala 30:58]
  assign _T_88 = _T_26 ? 22'h0 : ~_T_86; // @[primitives.scala 74:21]
  assign _T_90 = {~_T_88,3'h7}; // @[Cat.scala 30:58]
  assign _T_100 = {_T_28[0],_T_28[1],_T_28[2]}; // @[Cat.scala 30:58]
  assign _T_101 = _T_26 ? _T_100 : 3'h0; // @[primitives.scala 61:24]
  assign _T_102 = _T_24 ? _T_90 : {{22'd0}, _T_101}; // @[primitives.scala 66:24]
  assign _T_103 = _T_22 ? _T_102 : 25'h0; // @[primitives.scala 61:24]
  assign _GEN_3 = {{24'd0}, doShiftSigDown1}; // @[RoundAnyRawFNToRecFN.scala 157:23]
  assign _T_104 = _T_103 | _GEN_3; // @[RoundAnyRawFNToRecFN.scala 157:23]
  assign _T_105 = {_T_104,2'h3}; // @[Cat.scala 30:58]
  assign _T_107 = {1'h0,_T_105[26:1]}; // @[Cat.scala 30:58]
  assign _T_109 = ~_T_107 & _T_105; // @[RoundAnyRawFNToRecFN.scala 161:46]
  assign _T_110 = io_in_sig & _T_109; // @[RoundAnyRawFNToRecFN.scala 162:40]
  assign _T_111 = _T_110 != 27'h0; // @[RoundAnyRawFNToRecFN.scala 162:56]
  assign _T_112 = io_in_sig & _T_107; // @[RoundAnyRawFNToRecFN.scala 163:42]
  assign _T_113 = _T_112 != 27'h0; // @[RoundAnyRawFNToRecFN.scala 163:62]
  assign _T_114 = _T_111 | _T_113; // @[RoundAnyRawFNToRecFN.scala 164:36]
  assign _T_115 = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38]
  assign _T_116 = _T_115 & _T_111; // @[RoundAnyRawFNToRecFN.scala 167:67]
  assign _T_117 = roundMagUp & _T_114; // @[RoundAnyRawFNToRecFN.scala 169:29]
  assign _T_118 = _T_116 | _T_117; // @[RoundAnyRawFNToRecFN.scala 168:31]
  assign _T_119 = io_in_sig | _T_105; // @[RoundAnyRawFNToRecFN.scala 172:32]
  assign _T_121 = _T_119[26:2] + 25'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  assign _T_122 = roundingMode_near_even & _T_111; // @[RoundAnyRawFNToRecFN.scala 173:49]
  assign _T_124 = _T_122 & ~_T_113; // @[RoundAnyRawFNToRecFN.scala 173:64]
  assign _T_126 = _T_124 ? _T_105[26:1] : 26'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  assign _T_128 = _T_121 & ~_T_126; // @[RoundAnyRawFNToRecFN.scala 172:61]
  assign _T_130 = io_in_sig & ~_T_105; // @[RoundAnyRawFNToRecFN.scala 178:30]
  assign _T_132 = roundingMode_odd & _T_114; // @[RoundAnyRawFNToRecFN.scala 179:42]
  assign _T_134 = _T_132 ? _T_109[26:1] : 26'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  assign _GEN_4 = {{1'd0}, _T_130[26:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_135 = _GEN_4 | _T_134; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_136 = _T_118 ? _T_128 : _T_135; // @[RoundAnyRawFNToRecFN.scala 171:16]
  assign _T_138 = {1'b0,$signed(_T_136[25:24])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  assign _GEN_5 = {{7{_T_138[2]}},_T_138}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign _T_139 = $signed(io_in_sExp) + $signed(_GEN_5); // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign common_expOut = _T_139[8:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  assign common_fractOut = doShiftSigDown1 ? _T_136[23:1] : _T_136[22:0]; // @[RoundAnyRawFNToRecFN.scala 187:16]
  assign _T_144 = _T_139[10:7]; // @[RoundAnyRawFNToRecFN.scala 194:30]
  assign common_overflow = $signed(_T_144) >= 4'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50]
  assign common_totalUnderflow = $signed(_T_139) < 11'sh6b; // @[RoundAnyRawFNToRecFN.scala 198:31]
  assign _T_149 = doShiftSigDown1 ? io_in_sig[2] : io_in_sig[1]; // @[RoundAnyRawFNToRecFN.scala 201:16]
  assign _T_151 = doShiftSigDown1 & io_in_sig[2]; // @[RoundAnyRawFNToRecFN.scala 203:30]
  assign _T_153 = io_in_sig[1:0] != 2'h0; // @[RoundAnyRawFNToRecFN.scala 203:70]
  assign _T_154 = _T_151 | _T_153; // @[RoundAnyRawFNToRecFN.scala 203:49]
  assign _T_156 = _T_115 & _T_149; // @[RoundAnyRawFNToRecFN.scala 205:67]
  assign _T_157 = roundMagUp & _T_154; // @[RoundAnyRawFNToRecFN.scala 207:29]
  assign _T_158 = _T_156 | _T_157; // @[RoundAnyRawFNToRecFN.scala 206:46]
  assign _T_161 = doShiftSigDown1 ? _T_136[25] : _T_136[24]; // @[RoundAnyRawFNToRecFN.scala 209:16]
  assign _T_162 = io_in_sExp[9:8]; // @[RoundAnyRawFNToRecFN.scala 218:48]
  assign _T_163 = $signed(_T_162) <= 2'sh0; // @[RoundAnyRawFNToRecFN.scala 218:62]
  assign _T_164 = _T_114 & _T_163; // @[RoundAnyRawFNToRecFN.scala 218:32]
  assign _T_167 = doShiftSigDown1 ? _T_105[3] : _T_105[2]; // @[RoundAnyRawFNToRecFN.scala 219:30]
  assign _T_168 = _T_164 & _T_167; // @[RoundAnyRawFNToRecFN.scala 218:74]
  assign _T_172 = doShiftSigDown1 ? _T_105[4] : _T_105[3]; // @[RoundAnyRawFNToRecFN.scala 221:39]
  assign _T_174 = io_detectTininess & ~_T_172; // @[RoundAnyRawFNToRecFN.scala 220:77]
  assign _T_175 = _T_174 & _T_161; // @[RoundAnyRawFNToRecFN.scala 224:38]
  assign _T_176 = _T_175 & _T_111; // @[RoundAnyRawFNToRecFN.scala 225:45]
  assign _T_177 = _T_176 & _T_158; // @[RoundAnyRawFNToRecFN.scala 225:60]
  assign _T_179 = _T_168 & ~_T_177; // @[RoundAnyRawFNToRecFN.scala 219:76]
  assign common_underflow = common_totalUnderflow | _T_179; // @[RoundAnyRawFNToRecFN.scala 215:40]
  assign common_inexact = common_totalUnderflow | _T_114; // @[RoundAnyRawFNToRecFN.scala 228:49]
  assign isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34]
  assign notNaN_isSpecialInfOut = io_infiniteExc | io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 234:49]
  assign _T_184 = ~isNaNOut & ~notNaN_isSpecialInfOut; // @[RoundAnyRawFNToRecFN.scala 235:33]
  assign commonCase = _T_184 & ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:61]
  assign overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  assign underflow = commonCase & common_underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  assign _T_186 = commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  assign inexact = overflow | _T_186; // @[RoundAnyRawFNToRecFN.scala 238:28]
  assign overflow_roundMagUp = _T_115 | roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  assign _T_188 = commonCase & common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 243:20]
  assign _T_189 = roundMagUp | roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 243:60]
  assign pegMinNonzeroMagOut = _T_188 & _T_189; // @[RoundAnyRawFNToRecFN.scala 243:45]
  assign pegMaxFiniteMagOut = overflow & ~overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 244:39]
  assign _T_191 = overflow & overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 246:45]
  assign notNaN_isInfOut = notNaN_isSpecialInfOut | _T_191; // @[RoundAnyRawFNToRecFN.scala 246:32]
  assign signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22]
  assign _T_192 = io_in_isZero | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 251:32]
  assign _T_193 = _T_192 ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign _T_195 = common_expOut & ~_T_193; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign _T_197 = pegMinNonzeroMagOut ? 9'h194 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 255:18]
  assign _T_199 = _T_195 & ~_T_197; // @[RoundAnyRawFNToRecFN.scala 254:17]
  assign _T_200 = pegMaxFiniteMagOut ? 9'h80 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 259:18]
  assign _T_202 = _T_199 & ~_T_200; // @[RoundAnyRawFNToRecFN.scala 258:17]
  assign _T_203 = notNaN_isInfOut ? 9'h40 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  assign _T_205 = _T_202 & ~_T_203; // @[RoundAnyRawFNToRecFN.scala 262:17]
  assign _T_206 = pegMinNonzeroMagOut ? 9'h6b : 9'h0; // @[RoundAnyRawFNToRecFN.scala 267:16]
  assign _T_207 = _T_205 | _T_206; // @[RoundAnyRawFNToRecFN.scala 266:18]
  assign _T_208 = pegMaxFiniteMagOut ? 9'h17f : 9'h0; // @[RoundAnyRawFNToRecFN.scala 271:16]
  assign _T_209 = _T_207 | _T_208; // @[RoundAnyRawFNToRecFN.scala 270:15]
  assign _T_210 = notNaN_isInfOut ? 9'h180 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  assign _T_211 = _T_209 | _T_210; // @[RoundAnyRawFNToRecFN.scala 274:15]
  assign _T_212 = isNaNOut ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 276:16]
  assign expOut = _T_211 | _T_212; // @[RoundAnyRawFNToRecFN.scala 275:77]
  assign _T_213 = isNaNOut | io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 278:22]
  assign _T_214 = _T_213 | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 278:38]
  assign _T_215 = isNaNOut ? 23'h400000 : 23'h0; // @[RoundAnyRawFNToRecFN.scala 279:16]
  assign _T_216 = _T_214 ? _T_215 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign _T_218 = pegMaxFiniteMagOut ? 23'h7fffff : 23'h0; // @[Bitwise.scala 72:12]
  assign fractOut = _T_216 | _T_218; // @[RoundAnyRawFNToRecFN.scala 281:11]
  assign _T_219 = {signOut,expOut}; // @[Cat.scala 30:58]
  assign _T_221 = {underflow,inexact}; // @[Cat.scala 30:58]
  assign _T_223 = {io_invalidExc,io_infiniteExc,overflow}; // @[Cat.scala 30:58]
  assign io_out = {_T_219,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
  assign io_exceptionFlags = {_T_223,_T_221}; // @[RoundAnyRawFNToRecFN.scala 285:23]
  assign RoundAnyRawFNToRecFN_5_covSum = 30'h0;
  assign io_covSum = RoundAnyRawFNToRecFN_5_covSum;
  assign metaAssert = 1'h0;
endmodule
module RoundAnyRawFNToRecFN_6(
  input         io_invalidExc,
  input         io_infiniteExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [12:0] io_in_sExp,
  input  [55:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire  _T_11; // @[RoundAnyRawFNToRecFN.scala 96:27]
  wire  _T_13; // @[RoundAnyRawFNToRecFN.scala 96:63]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42]
  wire  doShiftSigDown1; // @[RoundAnyRawFNToRecFN.scala 118:61]
  wire  _T_22; // @[primitives.scala 57:25]
  wire  _T_24; // @[primitives.scala 57:25]
  wire  _T_26; // @[primitives.scala 57:25]
  wire  _T_28; // @[primitives.scala 57:25]
  wire  _T_30; // @[primitives.scala 57:25]
  wire  _T_32; // @[primitives.scala 57:25]
  wire [5:0] _T_33; // @[primitives.scala 58:26]
  wire [64:0] _T_34; // @[primitives.scala 77:58]
  wire [31:0] _T_40; // @[Bitwise.scala 103:31]
  wire [31:0] _T_42; // @[Bitwise.scala 103:65]
  wire [31:0] _T_44; // @[Bitwise.scala 103:75]
  wire [31:0] _T_45; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_0; // @[Bitwise.scala 103:31]
  wire [31:0] _T_50; // @[Bitwise.scala 103:31]
  wire [31:0] _T_52; // @[Bitwise.scala 103:65]
  wire [31:0] _T_54; // @[Bitwise.scala 103:75]
  wire [31:0] _T_55; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_1; // @[Bitwise.scala 103:31]
  wire [31:0] _T_60; // @[Bitwise.scala 103:31]
  wire [31:0] _T_62; // @[Bitwise.scala 103:65]
  wire [31:0] _T_64; // @[Bitwise.scala 103:75]
  wire [31:0] _T_65; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_2; // @[Bitwise.scala 103:31]
  wire [31:0] _T_70; // @[Bitwise.scala 103:31]
  wire [31:0] _T_72; // @[Bitwise.scala 103:65]
  wire [31:0] _T_74; // @[Bitwise.scala 103:75]
  wire [31:0] _T_75; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_3; // @[Bitwise.scala 103:31]
  wire [31:0] _T_80; // @[Bitwise.scala 103:31]
  wire [31:0] _T_82; // @[Bitwise.scala 103:65]
  wire [31:0] _T_84; // @[Bitwise.scala 103:75]
  wire [31:0] _T_85; // @[Bitwise.scala 103:39]
  wire [15:0] _T_91; // @[Bitwise.scala 103:31]
  wire [15:0] _T_93; // @[Bitwise.scala 103:65]
  wire [15:0] _T_95; // @[Bitwise.scala 103:75]
  wire [15:0] _T_96; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_4; // @[Bitwise.scala 103:31]
  wire [15:0] _T_101; // @[Bitwise.scala 103:31]
  wire [15:0] _T_103; // @[Bitwise.scala 103:65]
  wire [15:0] _T_105; // @[Bitwise.scala 103:75]
  wire [15:0] _T_106; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_5; // @[Bitwise.scala 103:31]
  wire [15:0] _T_111; // @[Bitwise.scala 103:31]
  wire [15:0] _T_113; // @[Bitwise.scala 103:65]
  wire [15:0] _T_115; // @[Bitwise.scala 103:75]
  wire [15:0] _T_116; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_6; // @[Bitwise.scala 103:31]
  wire [15:0] _T_121; // @[Bitwise.scala 103:31]
  wire [15:0] _T_123; // @[Bitwise.scala 103:65]
  wire [15:0] _T_125; // @[Bitwise.scala 103:75]
  wire [15:0] _T_126; // @[Bitwise.scala 103:39]
  wire [50:0] _T_135; // @[Cat.scala 30:58]
  wire [50:0] _T_137; // @[primitives.scala 74:21]
  wire [50:0] _T_140; // @[primitives.scala 74:21]
  wire [50:0] _T_143; // @[primitives.scala 74:21]
  wire [50:0] _T_146; // @[primitives.scala 74:21]
  wire [53:0] _T_148; // @[Cat.scala 30:58]
  wire [2:0] _T_164; // @[Cat.scala 30:58]
  wire [2:0] _T_165; // @[primitives.scala 61:24]
  wire [2:0] _T_166; // @[primitives.scala 61:24]
  wire [2:0] _T_167; // @[primitives.scala 61:24]
  wire [2:0] _T_168; // @[primitives.scala 61:24]
  wire [53:0] _T_169; // @[primitives.scala 66:24]
  wire [53:0] _T_170; // @[primitives.scala 61:24]
  wire [53:0] _GEN_7; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [53:0] _T_171; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [55:0] _T_172; // @[Cat.scala 30:58]
  wire [55:0] _T_174; // @[Cat.scala 30:58]
  wire [55:0] _T_176; // @[RoundAnyRawFNToRecFN.scala 161:46]
  wire [55:0] _T_177; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  _T_178; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [55:0] _T_179; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  _T_180; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  _T_181; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire  _T_182; // @[RoundAnyRawFNToRecFN.scala 167:38]
  wire  _T_183; // @[RoundAnyRawFNToRecFN.scala 167:67]
  wire  _T_184; // @[RoundAnyRawFNToRecFN.scala 169:29]
  wire  _T_185; // @[RoundAnyRawFNToRecFN.scala 168:31]
  wire [55:0] _T_186; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [54:0] _T_188; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _T_189; // @[RoundAnyRawFNToRecFN.scala 173:49]
  wire  _T_191; // @[RoundAnyRawFNToRecFN.scala 173:64]
  wire [54:0] _T_193; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [54:0] _T_195; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [55:0] _T_197; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire  _T_199; // @[RoundAnyRawFNToRecFN.scala 179:42]
  wire [54:0] _T_201; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [54:0] _GEN_8; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [54:0] _T_202; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [54:0] _T_203; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _T_205; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [12:0] _GEN_9; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [13:0] _T_206; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [11:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [51:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 187:16]
  wire [3:0] _T_211; // @[RoundAnyRawFNToRecFN.scala 194:30]
  wire  common_overflow; // @[RoundAnyRawFNToRecFN.scala 194:50]
  wire  common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 198:31]
  wire  _T_216; // @[RoundAnyRawFNToRecFN.scala 201:16]
  wire  _T_218; // @[RoundAnyRawFNToRecFN.scala 203:30]
  wire  _T_220; // @[RoundAnyRawFNToRecFN.scala 203:70]
  wire  _T_221; // @[RoundAnyRawFNToRecFN.scala 203:49]
  wire  _T_223; // @[RoundAnyRawFNToRecFN.scala 205:67]
  wire  _T_224; // @[RoundAnyRawFNToRecFN.scala 207:29]
  wire  _T_225; // @[RoundAnyRawFNToRecFN.scala 206:46]
  wire  _T_228; // @[RoundAnyRawFNToRecFN.scala 209:16]
  wire [1:0] _T_229; // @[RoundAnyRawFNToRecFN.scala 218:48]
  wire  _T_230; // @[RoundAnyRawFNToRecFN.scala 218:62]
  wire  _T_231; // @[RoundAnyRawFNToRecFN.scala 218:32]
  wire  _T_234; // @[RoundAnyRawFNToRecFN.scala 219:30]
  wire  _T_235; // @[RoundAnyRawFNToRecFN.scala 218:74]
  wire  _T_239; // @[RoundAnyRawFNToRecFN.scala 221:39]
  wire  _T_241; // @[RoundAnyRawFNToRecFN.scala 220:77]
  wire  _T_242; // @[RoundAnyRawFNToRecFN.scala 224:38]
  wire  _T_243; // @[RoundAnyRawFNToRecFN.scala 225:45]
  wire  _T_244; // @[RoundAnyRawFNToRecFN.scala 225:60]
  wire  _T_246; // @[RoundAnyRawFNToRecFN.scala 219:76]
  wire  common_underflow; // @[RoundAnyRawFNToRecFN.scala 215:40]
  wire  common_inexact; // @[RoundAnyRawFNToRecFN.scala 228:49]
  wire  isNaNOut; // @[RoundAnyRawFNToRecFN.scala 233:34]
  wire  notNaN_isSpecialInfOut; // @[RoundAnyRawFNToRecFN.scala 234:49]
  wire  _T_251; // @[RoundAnyRawFNToRecFN.scala 235:33]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:61]
  wire  overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  wire  underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  wire  _T_253; // @[RoundAnyRawFNToRecFN.scala 238:43]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:28]
  wire  overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  wire  _T_255; // @[RoundAnyRawFNToRecFN.scala 243:20]
  wire  _T_256; // @[RoundAnyRawFNToRecFN.scala 243:60]
  wire  pegMinNonzeroMagOut; // @[RoundAnyRawFNToRecFN.scala 243:45]
  wire  pegMaxFiniteMagOut; // @[RoundAnyRawFNToRecFN.scala 244:39]
  wire  _T_258; // @[RoundAnyRawFNToRecFN.scala 246:45]
  wire  notNaN_isInfOut; // @[RoundAnyRawFNToRecFN.scala 246:32]
  wire  signOut; // @[RoundAnyRawFNToRecFN.scala 248:22]
  wire  _T_259; // @[RoundAnyRawFNToRecFN.scala 251:32]
  wire [11:0] _T_260; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [11:0] _T_262; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [11:0] _T_264; // @[RoundAnyRawFNToRecFN.scala 255:18]
  wire [11:0] _T_266; // @[RoundAnyRawFNToRecFN.scala 254:17]
  wire [11:0] _T_267; // @[RoundAnyRawFNToRecFN.scala 259:18]
  wire [11:0] _T_269; // @[RoundAnyRawFNToRecFN.scala 258:17]
  wire [11:0] _T_270; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [11:0] _T_272; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [11:0] _T_273; // @[RoundAnyRawFNToRecFN.scala 267:16]
  wire [11:0] _T_274; // @[RoundAnyRawFNToRecFN.scala 266:18]
  wire [11:0] _T_275; // @[RoundAnyRawFNToRecFN.scala 271:16]
  wire [11:0] _T_276; // @[RoundAnyRawFNToRecFN.scala 270:15]
  wire [11:0] _T_277; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [11:0] _T_278; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [11:0] _T_279; // @[RoundAnyRawFNToRecFN.scala 276:16]
  wire [11:0] expOut; // @[RoundAnyRawFNToRecFN.scala 275:77]
  wire  _T_280; // @[RoundAnyRawFNToRecFN.scala 278:22]
  wire  _T_281; // @[RoundAnyRawFNToRecFN.scala 278:38]
  wire [51:0] _T_282; // @[RoundAnyRawFNToRecFN.scala 279:16]
  wire [51:0] _T_283; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [51:0] _T_285; // @[Bitwise.scala 72:12]
  wire [51:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 281:11]
  wire [12:0] _T_286; // @[Cat.scala 30:58]
  wire [1:0] _T_288; // @[Cat.scala 30:58]
  wire [2:0] _T_290; // @[Cat.scala 30:58]
  wire [29:0] RoundAnyRawFNToRecFN_6_covSum;
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53]
  assign roundingMode_odd = io_roundingMode == 3'h5; // @[RoundAnyRawFNToRecFN.scala 93:53]
  assign _T_11 = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27]
  assign _T_13 = roundingMode_max & ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:63]
  assign roundMagUp = _T_11 | _T_13; // @[RoundAnyRawFNToRecFN.scala 96:42]
  assign doShiftSigDown1 = io_in_sig[55]; // @[RoundAnyRawFNToRecFN.scala 118:61]
  assign _T_22 = ~io_in_sExp[11]; // @[primitives.scala 57:25]
  assign _T_24 = ~io_in_sExp[10]; // @[primitives.scala 57:25]
  assign _T_26 = ~io_in_sExp[9]; // @[primitives.scala 57:25]
  assign _T_28 = ~io_in_sExp[8]; // @[primitives.scala 57:25]
  assign _T_30 = ~io_in_sExp[7]; // @[primitives.scala 57:25]
  assign _T_32 = ~io_in_sExp[6]; // @[primitives.scala 57:25]
  assign _T_33 = ~io_in_sExp[5:0]; // @[primitives.scala 58:26]
  assign _T_34 = -65'sh10000000000000000 >>> _T_33; // @[primitives.scala 77:58]
  assign _T_40 = {{16'd0}, _T_34[44:29]}; // @[Bitwise.scala 103:31]
  assign _T_42 = {_T_34[28:13], 16'h0}; // @[Bitwise.scala 103:65]
  assign _T_44 = _T_42 & 32'hffff0000; // @[Bitwise.scala 103:75]
  assign _T_45 = _T_40 | _T_44; // @[Bitwise.scala 103:39]
  assign _GEN_0 = {{8'd0}, _T_45[31:8]}; // @[Bitwise.scala 103:31]
  assign _T_50 = _GEN_0 & 32'hff00ff; // @[Bitwise.scala 103:31]
  assign _T_52 = {_T_45[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_54 = _T_52 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  assign _T_55 = _T_50 | _T_54; // @[Bitwise.scala 103:39]
  assign _GEN_1 = {{4'd0}, _T_55[31:4]}; // @[Bitwise.scala 103:31]
  assign _T_60 = _GEN_1 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  assign _T_62 = {_T_55[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_64 = _T_62 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  assign _T_65 = _T_60 | _T_64; // @[Bitwise.scala 103:39]
  assign _GEN_2 = {{2'd0}, _T_65[31:2]}; // @[Bitwise.scala 103:31]
  assign _T_70 = _GEN_2 & 32'h33333333; // @[Bitwise.scala 103:31]
  assign _T_72 = {_T_65[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_74 = _T_72 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  assign _T_75 = _T_70 | _T_74; // @[Bitwise.scala 103:39]
  assign _GEN_3 = {{1'd0}, _T_75[31:1]}; // @[Bitwise.scala 103:31]
  assign _T_80 = _GEN_3 & 32'h55555555; // @[Bitwise.scala 103:31]
  assign _T_82 = {_T_75[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_84 = _T_82 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  assign _T_85 = _T_80 | _T_84; // @[Bitwise.scala 103:39]
  assign _T_91 = {{8'd0}, _T_34[60:53]}; // @[Bitwise.scala 103:31]
  assign _T_93 = {_T_34[52:45], 8'h0}; // @[Bitwise.scala 103:65]
  assign _T_95 = _T_93 & 16'hff00; // @[Bitwise.scala 103:75]
  assign _T_96 = _T_91 | _T_95; // @[Bitwise.scala 103:39]
  assign _GEN_4 = {{4'd0}, _T_96[15:4]}; // @[Bitwise.scala 103:31]
  assign _T_101 = _GEN_4 & 16'hf0f; // @[Bitwise.scala 103:31]
  assign _T_103 = {_T_96[11:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _T_105 = _T_103 & 16'hf0f0; // @[Bitwise.scala 103:75]
  assign _T_106 = _T_101 | _T_105; // @[Bitwise.scala 103:39]
  assign _GEN_5 = {{2'd0}, _T_106[15:2]}; // @[Bitwise.scala 103:31]
  assign _T_111 = _GEN_5 & 16'h3333; // @[Bitwise.scala 103:31]
  assign _T_113 = {_T_106[13:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _T_115 = _T_113 & 16'hcccc; // @[Bitwise.scala 103:75]
  assign _T_116 = _T_111 | _T_115; // @[Bitwise.scala 103:39]
  assign _GEN_6 = {{1'd0}, _T_116[15:1]}; // @[Bitwise.scala 103:31]
  assign _T_121 = _GEN_6 & 16'h5555; // @[Bitwise.scala 103:31]
  assign _T_123 = {_T_116[14:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _T_125 = _T_123 & 16'haaaa; // @[Bitwise.scala 103:75]
  assign _T_126 = _T_121 | _T_125; // @[Bitwise.scala 103:39]
  assign _T_135 = {_T_85,_T_126,_T_34[61],_T_34[62],_T_34[63]}; // @[Cat.scala 30:58]
  assign _T_137 = _T_32 ? 51'h0 : ~_T_135; // @[primitives.scala 74:21]
  assign _T_140 = _T_30 ? 51'h0 : _T_137[50:0]; // @[primitives.scala 74:21]
  assign _T_143 = _T_28 ? 51'h0 : _T_140[50:0]; // @[primitives.scala 74:21]
  assign _T_146 = _T_26 ? 51'h0 : _T_143[50:0]; // @[primitives.scala 74:21]
  assign _T_148 = {~_T_146,3'h7}; // @[Cat.scala 30:58]
  assign _T_164 = {_T_34[0],_T_34[1],_T_34[2]}; // @[Cat.scala 30:58]
  assign _T_165 = _T_32 ? _T_164 : 3'h0; // @[primitives.scala 61:24]
  assign _T_166 = _T_30 ? _T_165 : 3'h0; // @[primitives.scala 61:24]
  assign _T_167 = _T_28 ? _T_166 : 3'h0; // @[primitives.scala 61:24]
  assign _T_168 = _T_26 ? _T_167 : 3'h0; // @[primitives.scala 61:24]
  assign _T_169 = _T_24 ? _T_148 : {{51'd0}, _T_168}; // @[primitives.scala 66:24]
  assign _T_170 = _T_22 ? _T_169 : 54'h0; // @[primitives.scala 61:24]
  assign _GEN_7 = {{53'd0}, doShiftSigDown1}; // @[RoundAnyRawFNToRecFN.scala 157:23]
  assign _T_171 = _T_170 | _GEN_7; // @[RoundAnyRawFNToRecFN.scala 157:23]
  assign _T_172 = {_T_171,2'h3}; // @[Cat.scala 30:58]
  assign _T_174 = {1'h0,_T_172[55:1]}; // @[Cat.scala 30:58]
  assign _T_176 = ~_T_174 & _T_172; // @[RoundAnyRawFNToRecFN.scala 161:46]
  assign _T_177 = io_in_sig & _T_176; // @[RoundAnyRawFNToRecFN.scala 162:40]
  assign _T_178 = _T_177 != 56'h0; // @[RoundAnyRawFNToRecFN.scala 162:56]
  assign _T_179 = io_in_sig & _T_174; // @[RoundAnyRawFNToRecFN.scala 163:42]
  assign _T_180 = _T_179 != 56'h0; // @[RoundAnyRawFNToRecFN.scala 163:62]
  assign _T_181 = _T_178 | _T_180; // @[RoundAnyRawFNToRecFN.scala 164:36]
  assign _T_182 = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38]
  assign _T_183 = _T_182 & _T_178; // @[RoundAnyRawFNToRecFN.scala 167:67]
  assign _T_184 = roundMagUp & _T_181; // @[RoundAnyRawFNToRecFN.scala 169:29]
  assign _T_185 = _T_183 | _T_184; // @[RoundAnyRawFNToRecFN.scala 168:31]
  assign _T_186 = io_in_sig | _T_172; // @[RoundAnyRawFNToRecFN.scala 172:32]
  assign _T_188 = _T_186[55:2] + 54'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  assign _T_189 = roundingMode_near_even & _T_178; // @[RoundAnyRawFNToRecFN.scala 173:49]
  assign _T_191 = _T_189 & ~_T_180; // @[RoundAnyRawFNToRecFN.scala 173:64]
  assign _T_193 = _T_191 ? _T_172[55:1] : 55'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  assign _T_195 = _T_188 & ~_T_193; // @[RoundAnyRawFNToRecFN.scala 172:61]
  assign _T_197 = io_in_sig & ~_T_172; // @[RoundAnyRawFNToRecFN.scala 178:30]
  assign _T_199 = roundingMode_odd & _T_181; // @[RoundAnyRawFNToRecFN.scala 179:42]
  assign _T_201 = _T_199 ? _T_176[55:1] : 55'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  assign _GEN_8 = {{1'd0}, _T_197[55:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_202 = _GEN_8 | _T_201; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_203 = _T_185 ? _T_195 : _T_202; // @[RoundAnyRawFNToRecFN.scala 171:16]
  assign _T_205 = {1'b0,$signed(_T_203[54:53])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  assign _GEN_9 = {{10{_T_205[2]}},_T_205}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign _T_206 = $signed(io_in_sExp) + $signed(_GEN_9); // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign common_expOut = _T_206[11:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  assign common_fractOut = doShiftSigDown1 ? _T_203[52:1] : _T_203[51:0]; // @[RoundAnyRawFNToRecFN.scala 187:16]
  assign _T_211 = _T_206[13:10]; // @[RoundAnyRawFNToRecFN.scala 194:30]
  assign common_overflow = $signed(_T_211) >= 4'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50]
  assign common_totalUnderflow = $signed(_T_206) < 14'sh3ce; // @[RoundAnyRawFNToRecFN.scala 198:31]
  assign _T_216 = doShiftSigDown1 ? io_in_sig[2] : io_in_sig[1]; // @[RoundAnyRawFNToRecFN.scala 201:16]
  assign _T_218 = doShiftSigDown1 & io_in_sig[2]; // @[RoundAnyRawFNToRecFN.scala 203:30]
  assign _T_220 = io_in_sig[1:0] != 2'h0; // @[RoundAnyRawFNToRecFN.scala 203:70]
  assign _T_221 = _T_218 | _T_220; // @[RoundAnyRawFNToRecFN.scala 203:49]
  assign _T_223 = _T_182 & _T_216; // @[RoundAnyRawFNToRecFN.scala 205:67]
  assign _T_224 = roundMagUp & _T_221; // @[RoundAnyRawFNToRecFN.scala 207:29]
  assign _T_225 = _T_223 | _T_224; // @[RoundAnyRawFNToRecFN.scala 206:46]
  assign _T_228 = doShiftSigDown1 ? _T_203[54] : _T_203[53]; // @[RoundAnyRawFNToRecFN.scala 209:16]
  assign _T_229 = io_in_sExp[12:11]; // @[RoundAnyRawFNToRecFN.scala 218:48]
  assign _T_230 = $signed(_T_229) <= 2'sh0; // @[RoundAnyRawFNToRecFN.scala 218:62]
  assign _T_231 = _T_181 & _T_230; // @[RoundAnyRawFNToRecFN.scala 218:32]
  assign _T_234 = doShiftSigDown1 ? _T_172[3] : _T_172[2]; // @[RoundAnyRawFNToRecFN.scala 219:30]
  assign _T_235 = _T_231 & _T_234; // @[RoundAnyRawFNToRecFN.scala 218:74]
  assign _T_239 = doShiftSigDown1 ? _T_172[4] : _T_172[3]; // @[RoundAnyRawFNToRecFN.scala 221:39]
  assign _T_241 = io_detectTininess & ~_T_239; // @[RoundAnyRawFNToRecFN.scala 220:77]
  assign _T_242 = _T_241 & _T_228; // @[RoundAnyRawFNToRecFN.scala 224:38]
  assign _T_243 = _T_242 & _T_178; // @[RoundAnyRawFNToRecFN.scala 225:45]
  assign _T_244 = _T_243 & _T_225; // @[RoundAnyRawFNToRecFN.scala 225:60]
  assign _T_246 = _T_235 & ~_T_244; // @[RoundAnyRawFNToRecFN.scala 219:76]
  assign common_underflow = common_totalUnderflow | _T_246; // @[RoundAnyRawFNToRecFN.scala 215:40]
  assign common_inexact = common_totalUnderflow | _T_181; // @[RoundAnyRawFNToRecFN.scala 228:49]
  assign isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34]
  assign notNaN_isSpecialInfOut = io_infiniteExc | io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 234:49]
  assign _T_251 = ~isNaNOut & ~notNaN_isSpecialInfOut; // @[RoundAnyRawFNToRecFN.scala 235:33]
  assign commonCase = _T_251 & ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:61]
  assign overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  assign underflow = commonCase & common_underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  assign _T_253 = commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  assign inexact = overflow | _T_253; // @[RoundAnyRawFNToRecFN.scala 238:28]
  assign overflow_roundMagUp = _T_182 | roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  assign _T_255 = commonCase & common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 243:20]
  assign _T_256 = roundMagUp | roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 243:60]
  assign pegMinNonzeroMagOut = _T_255 & _T_256; // @[RoundAnyRawFNToRecFN.scala 243:45]
  assign pegMaxFiniteMagOut = overflow & ~overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 244:39]
  assign _T_258 = overflow & overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 246:45]
  assign notNaN_isInfOut = notNaN_isSpecialInfOut | _T_258; // @[RoundAnyRawFNToRecFN.scala 246:32]
  assign signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22]
  assign _T_259 = io_in_isZero | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 251:32]
  assign _T_260 = _T_259 ? 12'he00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign _T_262 = common_expOut & ~_T_260; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign _T_264 = pegMinNonzeroMagOut ? 12'hc31 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 255:18]
  assign _T_266 = _T_262 & ~_T_264; // @[RoundAnyRawFNToRecFN.scala 254:17]
  assign _T_267 = pegMaxFiniteMagOut ? 12'h400 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 259:18]
  assign _T_269 = _T_266 & ~_T_267; // @[RoundAnyRawFNToRecFN.scala 258:17]
  assign _T_270 = notNaN_isInfOut ? 12'h200 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  assign _T_272 = _T_269 & ~_T_270; // @[RoundAnyRawFNToRecFN.scala 262:17]
  assign _T_273 = pegMinNonzeroMagOut ? 12'h3ce : 12'h0; // @[RoundAnyRawFNToRecFN.scala 267:16]
  assign _T_274 = _T_272 | _T_273; // @[RoundAnyRawFNToRecFN.scala 266:18]
  assign _T_275 = pegMaxFiniteMagOut ? 12'hbff : 12'h0; // @[RoundAnyRawFNToRecFN.scala 271:16]
  assign _T_276 = _T_274 | _T_275; // @[RoundAnyRawFNToRecFN.scala 270:15]
  assign _T_277 = notNaN_isInfOut ? 12'hc00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  assign _T_278 = _T_276 | _T_277; // @[RoundAnyRawFNToRecFN.scala 274:15]
  assign _T_279 = isNaNOut ? 12'he00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 276:16]
  assign expOut = _T_278 | _T_279; // @[RoundAnyRawFNToRecFN.scala 275:77]
  assign _T_280 = isNaNOut | io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 278:22]
  assign _T_281 = _T_280 | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 278:38]
  assign _T_282 = isNaNOut ? 52'h8000000000000 : 52'h0; // @[RoundAnyRawFNToRecFN.scala 279:16]
  assign _T_283 = _T_281 ? _T_282 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign _T_285 = pegMaxFiniteMagOut ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  assign fractOut = _T_283 | _T_285; // @[RoundAnyRawFNToRecFN.scala 281:11]
  assign _T_286 = {signOut,expOut}; // @[Cat.scala 30:58]
  assign _T_288 = {underflow,inexact}; // @[Cat.scala 30:58]
  assign _T_290 = {io_invalidExc,io_infiniteExc,overflow}; // @[Cat.scala 30:58]
  assign io_out = {_T_286,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
  assign io_exceptionFlags = {_T_290,_T_288}; // @[RoundAnyRawFNToRecFN.scala 285:23]
  assign RoundAnyRawFNToRecFN_6_covSum = 30'h0;
  assign io_covSum = RoundAnyRawFNToRecFN_6_covSum;
  assign metaAssert = 1'h0;
endmodule
